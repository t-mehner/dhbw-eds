--------------------------------------------------------------------------------
-- Company: 
-- Engineer:
--
-- Create Date:   08:51:40 10/22/2018
-- Design Name:   
-- Module Name:   /home/torben/Documents/DHBW/EDS/Projekte/hw_mul_pipelined/hw_mul_pipelined_tb.vhd
-- Project Name:  hw_mul_pipelined
-- Target Device:  
-- Tool versions:  
-- Description:   
-- 
-- VHDL Test Bench Created by ISE for module: hw_mul_pipelined
-- 
-- Dependencies:
-- 
-- Revision:
-- Revision 0.01 - File Created
-- Additional Comments:
--
-- Notes: 
-- This testbench has been automatically generated using types std_logic and
-- std_logic_vector for the ports of the unit under test.  Xilinx recommends
-- that these types always be used for the top-level I/O of a design in order
-- to guarantee that the testbench will bind correctly to the post-implementation 
-- simulation model.
--------------------------------------------------------------------------------
LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
 
-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
USE ieee.numeric_std.ALL;
 
ENTITY hw_mul_pipelined_tb IS
END hw_mul_pipelined_tb;
 
ARCHITECTURE behavior OF hw_mul_pipelined_tb IS 
 
   -- Component Declaration for the Unit Under Test (UUT)    

   --Inputs
   signal reset : std_logic := '0';
   signal clk : std_logic := '0';
   signal valid_in : std_logic := '0';
   signal a : unsigned(7 downto 0) := (others => '0');
   signal b : unsigned(7 downto 0) := (others => '0');

 	--Outputs
   signal valid_out : std_logic;
   signal q : unsigned(15 downto 0);

   -- Clock period definitions
   constant clk_period : time := 10 ns;
 
	signal counter : integer := 0;
	
	type result_type is array (0 to 65535) of integer;
	
	constant results : result_type := (
		0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
0, 1, 2, 3, 4, 5, 6, 7, 8, 9, 10, 11, 12, 13, 14, 15, 16, 17, 18, 19, 20, 21, 22, 23, 24, 25, 26, 27, 28, 29, 30, 31, 32, 33, 34, 35, 36, 37, 38, 39, 40, 41, 42, 43, 44, 45, 46, 47, 48, 49, 50, 51, 52, 53, 54, 55, 56, 57, 58, 59, 60, 61, 62, 63, 64, 65, 66, 67, 68, 69, 70, 71, 72, 73, 74, 75, 76, 77, 78, 79, 80, 81, 82, 83, 84, 85, 86, 87, 88, 89, 90, 91, 92, 93, 94, 95, 96, 97, 98, 99, 100, 101, 102, 103, 104, 105, 106, 107, 108, 109, 110, 111, 112, 113, 114, 115, 116, 117, 118, 119, 120, 121, 122, 123, 124, 125, 126, 127, 128, 129, 130, 131, 132, 133, 134, 135, 136, 137, 138, 139, 140, 141, 142, 143, 144, 145, 146, 147, 148, 149, 150, 151, 152, 153, 154, 155, 156, 157, 158, 159, 160, 161, 162, 163, 164, 165, 166, 167, 168, 169, 170, 171, 172, 173, 174, 175, 176, 177, 178, 179, 180, 181, 182, 183, 184, 185, 186, 187, 188, 189, 190, 191, 192, 193, 194, 195, 196, 197, 198, 199, 200, 201, 202, 203, 204, 205, 206, 207, 208, 209, 210, 211, 212, 213, 214, 215, 216, 217, 218, 219, 220, 221, 222, 223, 224, 225, 226, 227, 228, 229, 230, 231, 232, 233, 234, 235, 236, 237, 238, 239, 240, 241, 242, 243, 244, 245, 246, 247, 248, 249, 250, 251, 252, 253, 254, 255, 
0, 2, 4, 6, 8, 10, 12, 14, 16, 18, 20, 22, 24, 26, 28, 30, 32, 34, 36, 38, 40, 42, 44, 46, 48, 50, 52, 54, 56, 58, 60, 62, 64, 66, 68, 70, 72, 74, 76, 78, 80, 82, 84, 86, 88, 90, 92, 94, 96, 98, 100, 102, 104, 106, 108, 110, 112, 114, 116, 118, 120, 122, 124, 126, 128, 130, 132, 134, 136, 138, 140, 142, 144, 146, 148, 150, 152, 154, 156, 158, 160, 162, 164, 166, 168, 170, 172, 174, 176, 178, 180, 182, 184, 186, 188, 190, 192, 194, 196, 198, 200, 202, 204, 206, 208, 210, 212, 214, 216, 218, 220, 222, 224, 226, 228, 230, 232, 234, 236, 238, 240, 242, 244, 246, 248, 250, 252, 254, 256, 258, 260, 262, 264, 266, 268, 270, 272, 274, 276, 278, 280, 282, 284, 286, 288, 290, 292, 294, 296, 298, 300, 302, 304, 306, 308, 310, 312, 314, 316, 318, 320, 322, 324, 326, 328, 330, 332, 334, 336, 338, 340, 342, 344, 346, 348, 350, 352, 354, 356, 358, 360, 362, 364, 366, 368, 370, 372, 374, 376, 378, 380, 382, 384, 386, 388, 390, 392, 394, 396, 398, 400, 402, 404, 406, 408, 410, 412, 414, 416, 418, 420, 422, 424, 426, 428, 430, 432, 434, 436, 438, 440, 442, 444, 446, 448, 450, 452, 454, 456, 458, 460, 462, 464, 466, 468, 470, 472, 474, 476, 478, 480, 482, 484, 486, 488, 490, 492, 494, 496, 498, 500, 502, 504, 506, 508, 510, 
0, 3, 6, 9, 12, 15, 18, 21, 24, 27, 30, 33, 36, 39, 42, 45, 48, 51, 54, 57, 60, 63, 66, 69, 72, 75, 78, 81, 84, 87, 90, 93, 96, 99, 102, 105, 108, 111, 114, 117, 120, 123, 126, 129, 132, 135, 138, 141, 144, 147, 150, 153, 156, 159, 162, 165, 168, 171, 174, 177, 180, 183, 186, 189, 192, 195, 198, 201, 204, 207, 210, 213, 216, 219, 222, 225, 228, 231, 234, 237, 240, 243, 246, 249, 252, 255, 258, 261, 264, 267, 270, 273, 276, 279, 282, 285, 288, 291, 294, 297, 300, 303, 306, 309, 312, 315, 318, 321, 324, 327, 330, 333, 336, 339, 342, 345, 348, 351, 354, 357, 360, 363, 366, 369, 372, 375, 378, 381, 384, 387, 390, 393, 396, 399, 402, 405, 408, 411, 414, 417, 420, 423, 426, 429, 432, 435, 438, 441, 444, 447, 450, 453, 456, 459, 462, 465, 468, 471, 474, 477, 480, 483, 486, 489, 492, 495, 498, 501, 504, 507, 510, 513, 516, 519, 522, 525, 528, 531, 534, 537, 540, 543, 546, 549, 552, 555, 558, 561, 564, 567, 570, 573, 576, 579, 582, 585, 588, 591, 594, 597, 600, 603, 606, 609, 612, 615, 618, 621, 624, 627, 630, 633, 636, 639, 642, 645, 648, 651, 654, 657, 660, 663, 666, 669, 672, 675, 678, 681, 684, 687, 690, 693, 696, 699, 702, 705, 708, 711, 714, 717, 720, 723, 726, 729, 732, 735, 738, 741, 744, 747, 750, 753, 756, 759, 762, 765, 
0, 4, 8, 12, 16, 20, 24, 28, 32, 36, 40, 44, 48, 52, 56, 60, 64, 68, 72, 76, 80, 84, 88, 92, 96, 100, 104, 108, 112, 116, 120, 124, 128, 132, 136, 140, 144, 148, 152, 156, 160, 164, 168, 172, 176, 180, 184, 188, 192, 196, 200, 204, 208, 212, 216, 220, 224, 228, 232, 236, 240, 244, 248, 252, 256, 260, 264, 268, 272, 276, 280, 284, 288, 292, 296, 300, 304, 308, 312, 316, 320, 324, 328, 332, 336, 340, 344, 348, 352, 356, 360, 364, 368, 372, 376, 380, 384, 388, 392, 396, 400, 404, 408, 412, 416, 420, 424, 428, 432, 436, 440, 444, 448, 452, 456, 460, 464, 468, 472, 476, 480, 484, 488, 492, 496, 500, 504, 508, 512, 516, 520, 524, 528, 532, 536, 540, 544, 548, 552, 556, 560, 564, 568, 572, 576, 580, 584, 588, 592, 596, 600, 604, 608, 612, 616, 620, 624, 628, 632, 636, 640, 644, 648, 652, 656, 660, 664, 668, 672, 676, 680, 684, 688, 692, 696, 700, 704, 708, 712, 716, 720, 724, 728, 732, 736, 740, 744, 748, 752, 756, 760, 764, 768, 772, 776, 780, 784, 788, 792, 796, 800, 804, 808, 812, 816, 820, 824, 828, 832, 836, 840, 844, 848, 852, 856, 860, 864, 868, 872, 876, 880, 884, 888, 892, 896, 900, 904, 908, 912, 916, 920, 924, 928, 932, 936, 940, 944, 948, 952, 956, 960, 964, 968, 972, 976, 980, 984, 988, 992, 996, 1000, 1004, 1008, 1012, 1016, 1020, 
0, 5, 10, 15, 20, 25, 30, 35, 40, 45, 50, 55, 60, 65, 70, 75, 80, 85, 90, 95, 100, 105, 110, 115, 120, 125, 130, 135, 140, 145, 150, 155, 160, 165, 170, 175, 180, 185, 190, 195, 200, 205, 210, 215, 220, 225, 230, 235, 240, 245, 250, 255, 260, 265, 270, 275, 280, 285, 290, 295, 300, 305, 310, 315, 320, 325, 330, 335, 340, 345, 350, 355, 360, 365, 370, 375, 380, 385, 390, 395, 400, 405, 410, 415, 420, 425, 430, 435, 440, 445, 450, 455, 460, 465, 470, 475, 480, 485, 490, 495, 500, 505, 510, 515, 520, 525, 530, 535, 540, 545, 550, 555, 560, 565, 570, 575, 580, 585, 590, 595, 600, 605, 610, 615, 620, 625, 630, 635, 640, 645, 650, 655, 660, 665, 670, 675, 680, 685, 690, 695, 700, 705, 710, 715, 720, 725, 730, 735, 740, 745, 750, 755, 760, 765, 770, 775, 780, 785, 790, 795, 800, 805, 810, 815, 820, 825, 830, 835, 840, 845, 850, 855, 860, 865, 870, 875, 880, 885, 890, 895, 900, 905, 910, 915, 920, 925, 930, 935, 940, 945, 950, 955, 960, 965, 970, 975, 980, 985, 990, 995, 1000, 1005, 1010, 1015, 1020, 1025, 1030, 1035, 1040, 1045, 1050, 1055, 1060, 1065, 1070, 1075, 1080, 1085, 1090, 1095, 1100, 1105, 1110, 1115, 1120, 1125, 1130, 1135, 1140, 1145, 1150, 1155, 1160, 1165, 1170, 1175, 1180, 1185, 1190, 1195, 1200, 1205, 1210, 1215, 1220, 1225, 1230, 1235, 1240, 1245, 1250, 1255, 1260, 1265, 1270, 1275, 
0, 6, 12, 18, 24, 30, 36, 42, 48, 54, 60, 66, 72, 78, 84, 90, 96, 102, 108, 114, 120, 126, 132, 138, 144, 150, 156, 162, 168, 174, 180, 186, 192, 198, 204, 210, 216, 222, 228, 234, 240, 246, 252, 258, 264, 270, 276, 282, 288, 294, 300, 306, 312, 318, 324, 330, 336, 342, 348, 354, 360, 366, 372, 378, 384, 390, 396, 402, 408, 414, 420, 426, 432, 438, 444, 450, 456, 462, 468, 474, 480, 486, 492, 498, 504, 510, 516, 522, 528, 534, 540, 546, 552, 558, 564, 570, 576, 582, 588, 594, 600, 606, 612, 618, 624, 630, 636, 642, 648, 654, 660, 666, 672, 678, 684, 690, 696, 702, 708, 714, 720, 726, 732, 738, 744, 750, 756, 762, 768, 774, 780, 786, 792, 798, 804, 810, 816, 822, 828, 834, 840, 846, 852, 858, 864, 870, 876, 882, 888, 894, 900, 906, 912, 918, 924, 930, 936, 942, 948, 954, 960, 966, 972, 978, 984, 990, 996, 1002, 1008, 1014, 1020, 1026, 1032, 1038, 1044, 1050, 1056, 1062, 1068, 1074, 1080, 1086, 1092, 1098, 1104, 1110, 1116, 1122, 1128, 1134, 1140, 1146, 1152, 1158, 1164, 1170, 1176, 1182, 1188, 1194, 1200, 1206, 1212, 1218, 1224, 1230, 1236, 1242, 1248, 1254, 1260, 1266, 1272, 1278, 1284, 1290, 1296, 1302, 1308, 1314, 1320, 1326, 1332, 1338, 1344, 1350, 1356, 1362, 1368, 1374, 1380, 1386, 1392, 1398, 1404, 1410, 1416, 1422, 1428, 1434, 1440, 1446, 1452, 1458, 1464, 1470, 1476, 1482, 1488, 1494, 1500, 1506, 1512, 1518, 1524, 1530, 
0, 7, 14, 21, 28, 35, 42, 49, 56, 63, 70, 77, 84, 91, 98, 105, 112, 119, 126, 133, 140, 147, 154, 161, 168, 175, 182, 189, 196, 203, 210, 217, 224, 231, 238, 245, 252, 259, 266, 273, 280, 287, 294, 301, 308, 315, 322, 329, 336, 343, 350, 357, 364, 371, 378, 385, 392, 399, 406, 413, 420, 427, 434, 441, 448, 455, 462, 469, 476, 483, 490, 497, 504, 511, 518, 525, 532, 539, 546, 553, 560, 567, 574, 581, 588, 595, 602, 609, 616, 623, 630, 637, 644, 651, 658, 665, 672, 679, 686, 693, 700, 707, 714, 721, 728, 735, 742, 749, 756, 763, 770, 777, 784, 791, 798, 805, 812, 819, 826, 833, 840, 847, 854, 861, 868, 875, 882, 889, 896, 903, 910, 917, 924, 931, 938, 945, 952, 959, 966, 973, 980, 987, 994, 1001, 1008, 1015, 1022, 1029, 1036, 1043, 1050, 1057, 1064, 1071, 1078, 1085, 1092, 1099, 1106, 1113, 1120, 1127, 1134, 1141, 1148, 1155, 1162, 1169, 1176, 1183, 1190, 1197, 1204, 1211, 1218, 1225, 1232, 1239, 1246, 1253, 1260, 1267, 1274, 1281, 1288, 1295, 1302, 1309, 1316, 1323, 1330, 1337, 1344, 1351, 1358, 1365, 1372, 1379, 1386, 1393, 1400, 1407, 1414, 1421, 1428, 1435, 1442, 1449, 1456, 1463, 1470, 1477, 1484, 1491, 1498, 1505, 1512, 1519, 1526, 1533, 1540, 1547, 1554, 1561, 1568, 1575, 1582, 1589, 1596, 1603, 1610, 1617, 1624, 1631, 1638, 1645, 1652, 1659, 1666, 1673, 1680, 1687, 1694, 1701, 1708, 1715, 1722, 1729, 1736, 1743, 1750, 1757, 1764, 1771, 1778, 1785, 
0, 8, 16, 24, 32, 40, 48, 56, 64, 72, 80, 88, 96, 104, 112, 120, 128, 136, 144, 152, 160, 168, 176, 184, 192, 200, 208, 216, 224, 232, 240, 248, 256, 264, 272, 280, 288, 296, 304, 312, 320, 328, 336, 344, 352, 360, 368, 376, 384, 392, 400, 408, 416, 424, 432, 440, 448, 456, 464, 472, 480, 488, 496, 504, 512, 520, 528, 536, 544, 552, 560, 568, 576, 584, 592, 600, 608, 616, 624, 632, 640, 648, 656, 664, 672, 680, 688, 696, 704, 712, 720, 728, 736, 744, 752, 760, 768, 776, 784, 792, 800, 808, 816, 824, 832, 840, 848, 856, 864, 872, 880, 888, 896, 904, 912, 920, 928, 936, 944, 952, 960, 968, 976, 984, 992, 1000, 1008, 1016, 1024, 1032, 1040, 1048, 1056, 1064, 1072, 1080, 1088, 1096, 1104, 1112, 1120, 1128, 1136, 1144, 1152, 1160, 1168, 1176, 1184, 1192, 1200, 1208, 1216, 1224, 1232, 1240, 1248, 1256, 1264, 1272, 1280, 1288, 1296, 1304, 1312, 1320, 1328, 1336, 1344, 1352, 1360, 1368, 1376, 1384, 1392, 1400, 1408, 1416, 1424, 1432, 1440, 1448, 1456, 1464, 1472, 1480, 1488, 1496, 1504, 1512, 1520, 1528, 1536, 1544, 1552, 1560, 1568, 1576, 1584, 1592, 1600, 1608, 1616, 1624, 1632, 1640, 1648, 1656, 1664, 1672, 1680, 1688, 1696, 1704, 1712, 1720, 1728, 1736, 1744, 1752, 1760, 1768, 1776, 1784, 1792, 1800, 1808, 1816, 1824, 1832, 1840, 1848, 1856, 1864, 1872, 1880, 1888, 1896, 1904, 1912, 1920, 1928, 1936, 1944, 1952, 1960, 1968, 1976, 1984, 1992, 2000, 2008, 2016, 2024, 2032, 2040, 
0, 9, 18, 27, 36, 45, 54, 63, 72, 81, 90, 99, 108, 117, 126, 135, 144, 153, 162, 171, 180, 189, 198, 207, 216, 225, 234, 243, 252, 261, 270, 279, 288, 297, 306, 315, 324, 333, 342, 351, 360, 369, 378, 387, 396, 405, 414, 423, 432, 441, 450, 459, 468, 477, 486, 495, 504, 513, 522, 531, 540, 549, 558, 567, 576, 585, 594, 603, 612, 621, 630, 639, 648, 657, 666, 675, 684, 693, 702, 711, 720, 729, 738, 747, 756, 765, 774, 783, 792, 801, 810, 819, 828, 837, 846, 855, 864, 873, 882, 891, 900, 909, 918, 927, 936, 945, 954, 963, 972, 981, 990, 999, 1008, 1017, 1026, 1035, 1044, 1053, 1062, 1071, 1080, 1089, 1098, 1107, 1116, 1125, 1134, 1143, 1152, 1161, 1170, 1179, 1188, 1197, 1206, 1215, 1224, 1233, 1242, 1251, 1260, 1269, 1278, 1287, 1296, 1305, 1314, 1323, 1332, 1341, 1350, 1359, 1368, 1377, 1386, 1395, 1404, 1413, 1422, 1431, 1440, 1449, 1458, 1467, 1476, 1485, 1494, 1503, 1512, 1521, 1530, 1539, 1548, 1557, 1566, 1575, 1584, 1593, 1602, 1611, 1620, 1629, 1638, 1647, 1656, 1665, 1674, 1683, 1692, 1701, 1710, 1719, 1728, 1737, 1746, 1755, 1764, 1773, 1782, 1791, 1800, 1809, 1818, 1827, 1836, 1845, 1854, 1863, 1872, 1881, 1890, 1899, 1908, 1917, 1926, 1935, 1944, 1953, 1962, 1971, 1980, 1989, 1998, 2007, 2016, 2025, 2034, 2043, 2052, 2061, 2070, 2079, 2088, 2097, 2106, 2115, 2124, 2133, 2142, 2151, 2160, 2169, 2178, 2187, 2196, 2205, 2214, 2223, 2232, 2241, 2250, 2259, 2268, 2277, 2286, 2295, 
0, 10, 20, 30, 40, 50, 60, 70, 80, 90, 100, 110, 120, 130, 140, 150, 160, 170, 180, 190, 200, 210, 220, 230, 240, 250, 260, 270, 280, 290, 300, 310, 320, 330, 340, 350, 360, 370, 380, 390, 400, 410, 420, 430, 440, 450, 460, 470, 480, 490, 500, 510, 520, 530, 540, 550, 560, 570, 580, 590, 600, 610, 620, 630, 640, 650, 660, 670, 680, 690, 700, 710, 720, 730, 740, 750, 760, 770, 780, 790, 800, 810, 820, 830, 840, 850, 860, 870, 880, 890, 900, 910, 920, 930, 940, 950, 960, 970, 980, 990, 1000, 1010, 1020, 1030, 1040, 1050, 1060, 1070, 1080, 1090, 1100, 1110, 1120, 1130, 1140, 1150, 1160, 1170, 1180, 1190, 1200, 1210, 1220, 1230, 1240, 1250, 1260, 1270, 1280, 1290, 1300, 1310, 1320, 1330, 1340, 1350, 1360, 1370, 1380, 1390, 1400, 1410, 1420, 1430, 1440, 1450, 1460, 1470, 1480, 1490, 1500, 1510, 1520, 1530, 1540, 1550, 1560, 1570, 1580, 1590, 1600, 1610, 1620, 1630, 1640, 1650, 1660, 1670, 1680, 1690, 1700, 1710, 1720, 1730, 1740, 1750, 1760, 1770, 1780, 1790, 1800, 1810, 1820, 1830, 1840, 1850, 1860, 1870, 1880, 1890, 1900, 1910, 1920, 1930, 1940, 1950, 1960, 1970, 1980, 1990, 2000, 2010, 2020, 2030, 2040, 2050, 2060, 2070, 2080, 2090, 2100, 2110, 2120, 2130, 2140, 2150, 2160, 2170, 2180, 2190, 2200, 2210, 2220, 2230, 2240, 2250, 2260, 2270, 2280, 2290, 2300, 2310, 2320, 2330, 2340, 2350, 2360, 2370, 2380, 2390, 2400, 2410, 2420, 2430, 2440, 2450, 2460, 2470, 2480, 2490, 2500, 2510, 2520, 2530, 2540, 2550, 
0, 11, 22, 33, 44, 55, 66, 77, 88, 99, 110, 121, 132, 143, 154, 165, 176, 187, 198, 209, 220, 231, 242, 253, 264, 275, 286, 297, 308, 319, 330, 341, 352, 363, 374, 385, 396, 407, 418, 429, 440, 451, 462, 473, 484, 495, 506, 517, 528, 539, 550, 561, 572, 583, 594, 605, 616, 627, 638, 649, 660, 671, 682, 693, 704, 715, 726, 737, 748, 759, 770, 781, 792, 803, 814, 825, 836, 847, 858, 869, 880, 891, 902, 913, 924, 935, 946, 957, 968, 979, 990, 1001, 1012, 1023, 1034, 1045, 1056, 1067, 1078, 1089, 1100, 1111, 1122, 1133, 1144, 1155, 1166, 1177, 1188, 1199, 1210, 1221, 1232, 1243, 1254, 1265, 1276, 1287, 1298, 1309, 1320, 1331, 1342, 1353, 1364, 1375, 1386, 1397, 1408, 1419, 1430, 1441, 1452, 1463, 1474, 1485, 1496, 1507, 1518, 1529, 1540, 1551, 1562, 1573, 1584, 1595, 1606, 1617, 1628, 1639, 1650, 1661, 1672, 1683, 1694, 1705, 1716, 1727, 1738, 1749, 1760, 1771, 1782, 1793, 1804, 1815, 1826, 1837, 1848, 1859, 1870, 1881, 1892, 1903, 1914, 1925, 1936, 1947, 1958, 1969, 1980, 1991, 2002, 2013, 2024, 2035, 2046, 2057, 2068, 2079, 2090, 2101, 2112, 2123, 2134, 2145, 2156, 2167, 2178, 2189, 2200, 2211, 2222, 2233, 2244, 2255, 2266, 2277, 2288, 2299, 2310, 2321, 2332, 2343, 2354, 2365, 2376, 2387, 2398, 2409, 2420, 2431, 2442, 2453, 2464, 2475, 2486, 2497, 2508, 2519, 2530, 2541, 2552, 2563, 2574, 2585, 2596, 2607, 2618, 2629, 2640, 2651, 2662, 2673, 2684, 2695, 2706, 2717, 2728, 2739, 2750, 2761, 2772, 2783, 2794, 2805, 
0, 12, 24, 36, 48, 60, 72, 84, 96, 108, 120, 132, 144, 156, 168, 180, 192, 204, 216, 228, 240, 252, 264, 276, 288, 300, 312, 324, 336, 348, 360, 372, 384, 396, 408, 420, 432, 444, 456, 468, 480, 492, 504, 516, 528, 540, 552, 564, 576, 588, 600, 612, 624, 636, 648, 660, 672, 684, 696, 708, 720, 732, 744, 756, 768, 780, 792, 804, 816, 828, 840, 852, 864, 876, 888, 900, 912, 924, 936, 948, 960, 972, 984, 996, 1008, 1020, 1032, 1044, 1056, 1068, 1080, 1092, 1104, 1116, 1128, 1140, 1152, 1164, 1176, 1188, 1200, 1212, 1224, 1236, 1248, 1260, 1272, 1284, 1296, 1308, 1320, 1332, 1344, 1356, 1368, 1380, 1392, 1404, 1416, 1428, 1440, 1452, 1464, 1476, 1488, 1500, 1512, 1524, 1536, 1548, 1560, 1572, 1584, 1596, 1608, 1620, 1632, 1644, 1656, 1668, 1680, 1692, 1704, 1716, 1728, 1740, 1752, 1764, 1776, 1788, 1800, 1812, 1824, 1836, 1848, 1860, 1872, 1884, 1896, 1908, 1920, 1932, 1944, 1956, 1968, 1980, 1992, 2004, 2016, 2028, 2040, 2052, 2064, 2076, 2088, 2100, 2112, 2124, 2136, 2148, 2160, 2172, 2184, 2196, 2208, 2220, 2232, 2244, 2256, 2268, 2280, 2292, 2304, 2316, 2328, 2340, 2352, 2364, 2376, 2388, 2400, 2412, 2424, 2436, 2448, 2460, 2472, 2484, 2496, 2508, 2520, 2532, 2544, 2556, 2568, 2580, 2592, 2604, 2616, 2628, 2640, 2652, 2664, 2676, 2688, 2700, 2712, 2724, 2736, 2748, 2760, 2772, 2784, 2796, 2808, 2820, 2832, 2844, 2856, 2868, 2880, 2892, 2904, 2916, 2928, 2940, 2952, 2964, 2976, 2988, 3000, 3012, 3024, 3036, 3048, 3060, 
0, 13, 26, 39, 52, 65, 78, 91, 104, 117, 130, 143, 156, 169, 182, 195, 208, 221, 234, 247, 260, 273, 286, 299, 312, 325, 338, 351, 364, 377, 390, 403, 416, 429, 442, 455, 468, 481, 494, 507, 520, 533, 546, 559, 572, 585, 598, 611, 624, 637, 650, 663, 676, 689, 702, 715, 728, 741, 754, 767, 780, 793, 806, 819, 832, 845, 858, 871, 884, 897, 910, 923, 936, 949, 962, 975, 988, 1001, 1014, 1027, 1040, 1053, 1066, 1079, 1092, 1105, 1118, 1131, 1144, 1157, 1170, 1183, 1196, 1209, 1222, 1235, 1248, 1261, 1274, 1287, 1300, 1313, 1326, 1339, 1352, 1365, 1378, 1391, 1404, 1417, 1430, 1443, 1456, 1469, 1482, 1495, 1508, 1521, 1534, 1547, 1560, 1573, 1586, 1599, 1612, 1625, 1638, 1651, 1664, 1677, 1690, 1703, 1716, 1729, 1742, 1755, 1768, 1781, 1794, 1807, 1820, 1833, 1846, 1859, 1872, 1885, 1898, 1911, 1924, 1937, 1950, 1963, 1976, 1989, 2002, 2015, 2028, 2041, 2054, 2067, 2080, 2093, 2106, 2119, 2132, 2145, 2158, 2171, 2184, 2197, 2210, 2223, 2236, 2249, 2262, 2275, 2288, 2301, 2314, 2327, 2340, 2353, 2366, 2379, 2392, 2405, 2418, 2431, 2444, 2457, 2470, 2483, 2496, 2509, 2522, 2535, 2548, 2561, 2574, 2587, 2600, 2613, 2626, 2639, 2652, 2665, 2678, 2691, 2704, 2717, 2730, 2743, 2756, 2769, 2782, 2795, 2808, 2821, 2834, 2847, 2860, 2873, 2886, 2899, 2912, 2925, 2938, 2951, 2964, 2977, 2990, 3003, 3016, 3029, 3042, 3055, 3068, 3081, 3094, 3107, 3120, 3133, 3146, 3159, 3172, 3185, 3198, 3211, 3224, 3237, 3250, 3263, 3276, 3289, 3302, 3315, 
0, 14, 28, 42, 56, 70, 84, 98, 112, 126, 140, 154, 168, 182, 196, 210, 224, 238, 252, 266, 280, 294, 308, 322, 336, 350, 364, 378, 392, 406, 420, 434, 448, 462, 476, 490, 504, 518, 532, 546, 560, 574, 588, 602, 616, 630, 644, 658, 672, 686, 700, 714, 728, 742, 756, 770, 784, 798, 812, 826, 840, 854, 868, 882, 896, 910, 924, 938, 952, 966, 980, 994, 1008, 1022, 1036, 1050, 1064, 1078, 1092, 1106, 1120, 1134, 1148, 1162, 1176, 1190, 1204, 1218, 1232, 1246, 1260, 1274, 1288, 1302, 1316, 1330, 1344, 1358, 1372, 1386, 1400, 1414, 1428, 1442, 1456, 1470, 1484, 1498, 1512, 1526, 1540, 1554, 1568, 1582, 1596, 1610, 1624, 1638, 1652, 1666, 1680, 1694, 1708, 1722, 1736, 1750, 1764, 1778, 1792, 1806, 1820, 1834, 1848, 1862, 1876, 1890, 1904, 1918, 1932, 1946, 1960, 1974, 1988, 2002, 2016, 2030, 2044, 2058, 2072, 2086, 2100, 2114, 2128, 2142, 2156, 2170, 2184, 2198, 2212, 2226, 2240, 2254, 2268, 2282, 2296, 2310, 2324, 2338, 2352, 2366, 2380, 2394, 2408, 2422, 2436, 2450, 2464, 2478, 2492, 2506, 2520, 2534, 2548, 2562, 2576, 2590, 2604, 2618, 2632, 2646, 2660, 2674, 2688, 2702, 2716, 2730, 2744, 2758, 2772, 2786, 2800, 2814, 2828, 2842, 2856, 2870, 2884, 2898, 2912, 2926, 2940, 2954, 2968, 2982, 2996, 3010, 3024, 3038, 3052, 3066, 3080, 3094, 3108, 3122, 3136, 3150, 3164, 3178, 3192, 3206, 3220, 3234, 3248, 3262, 3276, 3290, 3304, 3318, 3332, 3346, 3360, 3374, 3388, 3402, 3416, 3430, 3444, 3458, 3472, 3486, 3500, 3514, 3528, 3542, 3556, 3570, 
0, 15, 30, 45, 60, 75, 90, 105, 120, 135, 150, 165, 180, 195, 210, 225, 240, 255, 270, 285, 300, 315, 330, 345, 360, 375, 390, 405, 420, 435, 450, 465, 480, 495, 510, 525, 540, 555, 570, 585, 600, 615, 630, 645, 660, 675, 690, 705, 720, 735, 750, 765, 780, 795, 810, 825, 840, 855, 870, 885, 900, 915, 930, 945, 960, 975, 990, 1005, 1020, 1035, 1050, 1065, 1080, 1095, 1110, 1125, 1140, 1155, 1170, 1185, 1200, 1215, 1230, 1245, 1260, 1275, 1290, 1305, 1320, 1335, 1350, 1365, 1380, 1395, 1410, 1425, 1440, 1455, 1470, 1485, 1500, 1515, 1530, 1545, 1560, 1575, 1590, 1605, 1620, 1635, 1650, 1665, 1680, 1695, 1710, 1725, 1740, 1755, 1770, 1785, 1800, 1815, 1830, 1845, 1860, 1875, 1890, 1905, 1920, 1935, 1950, 1965, 1980, 1995, 2010, 2025, 2040, 2055, 2070, 2085, 2100, 2115, 2130, 2145, 2160, 2175, 2190, 2205, 2220, 2235, 2250, 2265, 2280, 2295, 2310, 2325, 2340, 2355, 2370, 2385, 2400, 2415, 2430, 2445, 2460, 2475, 2490, 2505, 2520, 2535, 2550, 2565, 2580, 2595, 2610, 2625, 2640, 2655, 2670, 2685, 2700, 2715, 2730, 2745, 2760, 2775, 2790, 2805, 2820, 2835, 2850, 2865, 2880, 2895, 2910, 2925, 2940, 2955, 2970, 2985, 3000, 3015, 3030, 3045, 3060, 3075, 3090, 3105, 3120, 3135, 3150, 3165, 3180, 3195, 3210, 3225, 3240, 3255, 3270, 3285, 3300, 3315, 3330, 3345, 3360, 3375, 3390, 3405, 3420, 3435, 3450, 3465, 3480, 3495, 3510, 3525, 3540, 3555, 3570, 3585, 3600, 3615, 3630, 3645, 3660, 3675, 3690, 3705, 3720, 3735, 3750, 3765, 3780, 3795, 3810, 3825, 
0, 16, 32, 48, 64, 80, 96, 112, 128, 144, 160, 176, 192, 208, 224, 240, 256, 272, 288, 304, 320, 336, 352, 368, 384, 400, 416, 432, 448, 464, 480, 496, 512, 528, 544, 560, 576, 592, 608, 624, 640, 656, 672, 688, 704, 720, 736, 752, 768, 784, 800, 816, 832, 848, 864, 880, 896, 912, 928, 944, 960, 976, 992, 1008, 1024, 1040, 1056, 1072, 1088, 1104, 1120, 1136, 1152, 1168, 1184, 1200, 1216, 1232, 1248, 1264, 1280, 1296, 1312, 1328, 1344, 1360, 1376, 1392, 1408, 1424, 1440, 1456, 1472, 1488, 1504, 1520, 1536, 1552, 1568, 1584, 1600, 1616, 1632, 1648, 1664, 1680, 1696, 1712, 1728, 1744, 1760, 1776, 1792, 1808, 1824, 1840, 1856, 1872, 1888, 1904, 1920, 1936, 1952, 1968, 1984, 2000, 2016, 2032, 2048, 2064, 2080, 2096, 2112, 2128, 2144, 2160, 2176, 2192, 2208, 2224, 2240, 2256, 2272, 2288, 2304, 2320, 2336, 2352, 2368, 2384, 2400, 2416, 2432, 2448, 2464, 2480, 2496, 2512, 2528, 2544, 2560, 2576, 2592, 2608, 2624, 2640, 2656, 2672, 2688, 2704, 2720, 2736, 2752, 2768, 2784, 2800, 2816, 2832, 2848, 2864, 2880, 2896, 2912, 2928, 2944, 2960, 2976, 2992, 3008, 3024, 3040, 3056, 3072, 3088, 3104, 3120, 3136, 3152, 3168, 3184, 3200, 3216, 3232, 3248, 3264, 3280, 3296, 3312, 3328, 3344, 3360, 3376, 3392, 3408, 3424, 3440, 3456, 3472, 3488, 3504, 3520, 3536, 3552, 3568, 3584, 3600, 3616, 3632, 3648, 3664, 3680, 3696, 3712, 3728, 3744, 3760, 3776, 3792, 3808, 3824, 3840, 3856, 3872, 3888, 3904, 3920, 3936, 3952, 3968, 3984, 4000, 4016, 4032, 4048, 4064, 4080, 
0, 17, 34, 51, 68, 85, 102, 119, 136, 153, 170, 187, 204, 221, 238, 255, 272, 289, 306, 323, 340, 357, 374, 391, 408, 425, 442, 459, 476, 493, 510, 527, 544, 561, 578, 595, 612, 629, 646, 663, 680, 697, 714, 731, 748, 765, 782, 799, 816, 833, 850, 867, 884, 901, 918, 935, 952, 969, 986, 1003, 1020, 1037, 1054, 1071, 1088, 1105, 1122, 1139, 1156, 1173, 1190, 1207, 1224, 1241, 1258, 1275, 1292, 1309, 1326, 1343, 1360, 1377, 1394, 1411, 1428, 1445, 1462, 1479, 1496, 1513, 1530, 1547, 1564, 1581, 1598, 1615, 1632, 1649, 1666, 1683, 1700, 1717, 1734, 1751, 1768, 1785, 1802, 1819, 1836, 1853, 1870, 1887, 1904, 1921, 1938, 1955, 1972, 1989, 2006, 2023, 2040, 2057, 2074, 2091, 2108, 2125, 2142, 2159, 2176, 2193, 2210, 2227, 2244, 2261, 2278, 2295, 2312, 2329, 2346, 2363, 2380, 2397, 2414, 2431, 2448, 2465, 2482, 2499, 2516, 2533, 2550, 2567, 2584, 2601, 2618, 2635, 2652, 2669, 2686, 2703, 2720, 2737, 2754, 2771, 2788, 2805, 2822, 2839, 2856, 2873, 2890, 2907, 2924, 2941, 2958, 2975, 2992, 3009, 3026, 3043, 3060, 3077, 3094, 3111, 3128, 3145, 3162, 3179, 3196, 3213, 3230, 3247, 3264, 3281, 3298, 3315, 3332, 3349, 3366, 3383, 3400, 3417, 3434, 3451, 3468, 3485, 3502, 3519, 3536, 3553, 3570, 3587, 3604, 3621, 3638, 3655, 3672, 3689, 3706, 3723, 3740, 3757, 3774, 3791, 3808, 3825, 3842, 3859, 3876, 3893, 3910, 3927, 3944, 3961, 3978, 3995, 4012, 4029, 4046, 4063, 4080, 4097, 4114, 4131, 4148, 4165, 4182, 4199, 4216, 4233, 4250, 4267, 4284, 4301, 4318, 4335, 
0, 18, 36, 54, 72, 90, 108, 126, 144, 162, 180, 198, 216, 234, 252, 270, 288, 306, 324, 342, 360, 378, 396, 414, 432, 450, 468, 486, 504, 522, 540, 558, 576, 594, 612, 630, 648, 666, 684, 702, 720, 738, 756, 774, 792, 810, 828, 846, 864, 882, 900, 918, 936, 954, 972, 990, 1008, 1026, 1044, 1062, 1080, 1098, 1116, 1134, 1152, 1170, 1188, 1206, 1224, 1242, 1260, 1278, 1296, 1314, 1332, 1350, 1368, 1386, 1404, 1422, 1440, 1458, 1476, 1494, 1512, 1530, 1548, 1566, 1584, 1602, 1620, 1638, 1656, 1674, 1692, 1710, 1728, 1746, 1764, 1782, 1800, 1818, 1836, 1854, 1872, 1890, 1908, 1926, 1944, 1962, 1980, 1998, 2016, 2034, 2052, 2070, 2088, 2106, 2124, 2142, 2160, 2178, 2196, 2214, 2232, 2250, 2268, 2286, 2304, 2322, 2340, 2358, 2376, 2394, 2412, 2430, 2448, 2466, 2484, 2502, 2520, 2538, 2556, 2574, 2592, 2610, 2628, 2646, 2664, 2682, 2700, 2718, 2736, 2754, 2772, 2790, 2808, 2826, 2844, 2862, 2880, 2898, 2916, 2934, 2952, 2970, 2988, 3006, 3024, 3042, 3060, 3078, 3096, 3114, 3132, 3150, 3168, 3186, 3204, 3222, 3240, 3258, 3276, 3294, 3312, 3330, 3348, 3366, 3384, 3402, 3420, 3438, 3456, 3474, 3492, 3510, 3528, 3546, 3564, 3582, 3600, 3618, 3636, 3654, 3672, 3690, 3708, 3726, 3744, 3762, 3780, 3798, 3816, 3834, 3852, 3870, 3888, 3906, 3924, 3942, 3960, 3978, 3996, 4014, 4032, 4050, 4068, 4086, 4104, 4122, 4140, 4158, 4176, 4194, 4212, 4230, 4248, 4266, 4284, 4302, 4320, 4338, 4356, 4374, 4392, 4410, 4428, 4446, 4464, 4482, 4500, 4518, 4536, 4554, 4572, 4590, 
0, 19, 38, 57, 76, 95, 114, 133, 152, 171, 190, 209, 228, 247, 266, 285, 304, 323, 342, 361, 380, 399, 418, 437, 456, 475, 494, 513, 532, 551, 570, 589, 608, 627, 646, 665, 684, 703, 722, 741, 760, 779, 798, 817, 836, 855, 874, 893, 912, 931, 950, 969, 988, 1007, 1026, 1045, 1064, 1083, 1102, 1121, 1140, 1159, 1178, 1197, 1216, 1235, 1254, 1273, 1292, 1311, 1330, 1349, 1368, 1387, 1406, 1425, 1444, 1463, 1482, 1501, 1520, 1539, 1558, 1577, 1596, 1615, 1634, 1653, 1672, 1691, 1710, 1729, 1748, 1767, 1786, 1805, 1824, 1843, 1862, 1881, 1900, 1919, 1938, 1957, 1976, 1995, 2014, 2033, 2052, 2071, 2090, 2109, 2128, 2147, 2166, 2185, 2204, 2223, 2242, 2261, 2280, 2299, 2318, 2337, 2356, 2375, 2394, 2413, 2432, 2451, 2470, 2489, 2508, 2527, 2546, 2565, 2584, 2603, 2622, 2641, 2660, 2679, 2698, 2717, 2736, 2755, 2774, 2793, 2812, 2831, 2850, 2869, 2888, 2907, 2926, 2945, 2964, 2983, 3002, 3021, 3040, 3059, 3078, 3097, 3116, 3135, 3154, 3173, 3192, 3211, 3230, 3249, 3268, 3287, 3306, 3325, 3344, 3363, 3382, 3401, 3420, 3439, 3458, 3477, 3496, 3515, 3534, 3553, 3572, 3591, 3610, 3629, 3648, 3667, 3686, 3705, 3724, 3743, 3762, 3781, 3800, 3819, 3838, 3857, 3876, 3895, 3914, 3933, 3952, 3971, 3990, 4009, 4028, 4047, 4066, 4085, 4104, 4123, 4142, 4161, 4180, 4199, 4218, 4237, 4256, 4275, 4294, 4313, 4332, 4351, 4370, 4389, 4408, 4427, 4446, 4465, 4484, 4503, 4522, 4541, 4560, 4579, 4598, 4617, 4636, 4655, 4674, 4693, 4712, 4731, 4750, 4769, 4788, 4807, 4826, 4845, 
0, 20, 40, 60, 80, 100, 120, 140, 160, 180, 200, 220, 240, 260, 280, 300, 320, 340, 360, 380, 400, 420, 440, 460, 480, 500, 520, 540, 560, 580, 600, 620, 640, 660, 680, 700, 720, 740, 760, 780, 800, 820, 840, 860, 880, 900, 920, 940, 960, 980, 1000, 1020, 1040, 1060, 1080, 1100, 1120, 1140, 1160, 1180, 1200, 1220, 1240, 1260, 1280, 1300, 1320, 1340, 1360, 1380, 1400, 1420, 1440, 1460, 1480, 1500, 1520, 1540, 1560, 1580, 1600, 1620, 1640, 1660, 1680, 1700, 1720, 1740, 1760, 1780, 1800, 1820, 1840, 1860, 1880, 1900, 1920, 1940, 1960, 1980, 2000, 2020, 2040, 2060, 2080, 2100, 2120, 2140, 2160, 2180, 2200, 2220, 2240, 2260, 2280, 2300, 2320, 2340, 2360, 2380, 2400, 2420, 2440, 2460, 2480, 2500, 2520, 2540, 2560, 2580, 2600, 2620, 2640, 2660, 2680, 2700, 2720, 2740, 2760, 2780, 2800, 2820, 2840, 2860, 2880, 2900, 2920, 2940, 2960, 2980, 3000, 3020, 3040, 3060, 3080, 3100, 3120, 3140, 3160, 3180, 3200, 3220, 3240, 3260, 3280, 3300, 3320, 3340, 3360, 3380, 3400, 3420, 3440, 3460, 3480, 3500, 3520, 3540, 3560, 3580, 3600, 3620, 3640, 3660, 3680, 3700, 3720, 3740, 3760, 3780, 3800, 3820, 3840, 3860, 3880, 3900, 3920, 3940, 3960, 3980, 4000, 4020, 4040, 4060, 4080, 4100, 4120, 4140, 4160, 4180, 4200, 4220, 4240, 4260, 4280, 4300, 4320, 4340, 4360, 4380, 4400, 4420, 4440, 4460, 4480, 4500, 4520, 4540, 4560, 4580, 4600, 4620, 4640, 4660, 4680, 4700, 4720, 4740, 4760, 4780, 4800, 4820, 4840, 4860, 4880, 4900, 4920, 4940, 4960, 4980, 5000, 5020, 5040, 5060, 5080, 5100, 
0, 21, 42, 63, 84, 105, 126, 147, 168, 189, 210, 231, 252, 273, 294, 315, 336, 357, 378, 399, 420, 441, 462, 483, 504, 525, 546, 567, 588, 609, 630, 651, 672, 693, 714, 735, 756, 777, 798, 819, 840, 861, 882, 903, 924, 945, 966, 987, 1008, 1029, 1050, 1071, 1092, 1113, 1134, 1155, 1176, 1197, 1218, 1239, 1260, 1281, 1302, 1323, 1344, 1365, 1386, 1407, 1428, 1449, 1470, 1491, 1512, 1533, 1554, 1575, 1596, 1617, 1638, 1659, 1680, 1701, 1722, 1743, 1764, 1785, 1806, 1827, 1848, 1869, 1890, 1911, 1932, 1953, 1974, 1995, 2016, 2037, 2058, 2079, 2100, 2121, 2142, 2163, 2184, 2205, 2226, 2247, 2268, 2289, 2310, 2331, 2352, 2373, 2394, 2415, 2436, 2457, 2478, 2499, 2520, 2541, 2562, 2583, 2604, 2625, 2646, 2667, 2688, 2709, 2730, 2751, 2772, 2793, 2814, 2835, 2856, 2877, 2898, 2919, 2940, 2961, 2982, 3003, 3024, 3045, 3066, 3087, 3108, 3129, 3150, 3171, 3192, 3213, 3234, 3255, 3276, 3297, 3318, 3339, 3360, 3381, 3402, 3423, 3444, 3465, 3486, 3507, 3528, 3549, 3570, 3591, 3612, 3633, 3654, 3675, 3696, 3717, 3738, 3759, 3780, 3801, 3822, 3843, 3864, 3885, 3906, 3927, 3948, 3969, 3990, 4011, 4032, 4053, 4074, 4095, 4116, 4137, 4158, 4179, 4200, 4221, 4242, 4263, 4284, 4305, 4326, 4347, 4368, 4389, 4410, 4431, 4452, 4473, 4494, 4515, 4536, 4557, 4578, 4599, 4620, 4641, 4662, 4683, 4704, 4725, 4746, 4767, 4788, 4809, 4830, 4851, 4872, 4893, 4914, 4935, 4956, 4977, 4998, 5019, 5040, 5061, 5082, 5103, 5124, 5145, 5166, 5187, 5208, 5229, 5250, 5271, 5292, 5313, 5334, 5355, 
0, 22, 44, 66, 88, 110, 132, 154, 176, 198, 220, 242, 264, 286, 308, 330, 352, 374, 396, 418, 440, 462, 484, 506, 528, 550, 572, 594, 616, 638, 660, 682, 704, 726, 748, 770, 792, 814, 836, 858, 880, 902, 924, 946, 968, 990, 1012, 1034, 1056, 1078, 1100, 1122, 1144, 1166, 1188, 1210, 1232, 1254, 1276, 1298, 1320, 1342, 1364, 1386, 1408, 1430, 1452, 1474, 1496, 1518, 1540, 1562, 1584, 1606, 1628, 1650, 1672, 1694, 1716, 1738, 1760, 1782, 1804, 1826, 1848, 1870, 1892, 1914, 1936, 1958, 1980, 2002, 2024, 2046, 2068, 2090, 2112, 2134, 2156, 2178, 2200, 2222, 2244, 2266, 2288, 2310, 2332, 2354, 2376, 2398, 2420, 2442, 2464, 2486, 2508, 2530, 2552, 2574, 2596, 2618, 2640, 2662, 2684, 2706, 2728, 2750, 2772, 2794, 2816, 2838, 2860, 2882, 2904, 2926, 2948, 2970, 2992, 3014, 3036, 3058, 3080, 3102, 3124, 3146, 3168, 3190, 3212, 3234, 3256, 3278, 3300, 3322, 3344, 3366, 3388, 3410, 3432, 3454, 3476, 3498, 3520, 3542, 3564, 3586, 3608, 3630, 3652, 3674, 3696, 3718, 3740, 3762, 3784, 3806, 3828, 3850, 3872, 3894, 3916, 3938, 3960, 3982, 4004, 4026, 4048, 4070, 4092, 4114, 4136, 4158, 4180, 4202, 4224, 4246, 4268, 4290, 4312, 4334, 4356, 4378, 4400, 4422, 4444, 4466, 4488, 4510, 4532, 4554, 4576, 4598, 4620, 4642, 4664, 4686, 4708, 4730, 4752, 4774, 4796, 4818, 4840, 4862, 4884, 4906, 4928, 4950, 4972, 4994, 5016, 5038, 5060, 5082, 5104, 5126, 5148, 5170, 5192, 5214, 5236, 5258, 5280, 5302, 5324, 5346, 5368, 5390, 5412, 5434, 5456, 5478, 5500, 5522, 5544, 5566, 5588, 5610, 
0, 23, 46, 69, 92, 115, 138, 161, 184, 207, 230, 253, 276, 299, 322, 345, 368, 391, 414, 437, 460, 483, 506, 529, 552, 575, 598, 621, 644, 667, 690, 713, 736, 759, 782, 805, 828, 851, 874, 897, 920, 943, 966, 989, 1012, 1035, 1058, 1081, 1104, 1127, 1150, 1173, 1196, 1219, 1242, 1265, 1288, 1311, 1334, 1357, 1380, 1403, 1426, 1449, 1472, 1495, 1518, 1541, 1564, 1587, 1610, 1633, 1656, 1679, 1702, 1725, 1748, 1771, 1794, 1817, 1840, 1863, 1886, 1909, 1932, 1955, 1978, 2001, 2024, 2047, 2070, 2093, 2116, 2139, 2162, 2185, 2208, 2231, 2254, 2277, 2300, 2323, 2346, 2369, 2392, 2415, 2438, 2461, 2484, 2507, 2530, 2553, 2576, 2599, 2622, 2645, 2668, 2691, 2714, 2737, 2760, 2783, 2806, 2829, 2852, 2875, 2898, 2921, 2944, 2967, 2990, 3013, 3036, 3059, 3082, 3105, 3128, 3151, 3174, 3197, 3220, 3243, 3266, 3289, 3312, 3335, 3358, 3381, 3404, 3427, 3450, 3473, 3496, 3519, 3542, 3565, 3588, 3611, 3634, 3657, 3680, 3703, 3726, 3749, 3772, 3795, 3818, 3841, 3864, 3887, 3910, 3933, 3956, 3979, 4002, 4025, 4048, 4071, 4094, 4117, 4140, 4163, 4186, 4209, 4232, 4255, 4278, 4301, 4324, 4347, 4370, 4393, 4416, 4439, 4462, 4485, 4508, 4531, 4554, 4577, 4600, 4623, 4646, 4669, 4692, 4715, 4738, 4761, 4784, 4807, 4830, 4853, 4876, 4899, 4922, 4945, 4968, 4991, 5014, 5037, 5060, 5083, 5106, 5129, 5152, 5175, 5198, 5221, 5244, 5267, 5290, 5313, 5336, 5359, 5382, 5405, 5428, 5451, 5474, 5497, 5520, 5543, 5566, 5589, 5612, 5635, 5658, 5681, 5704, 5727, 5750, 5773, 5796, 5819, 5842, 5865, 
0, 24, 48, 72, 96, 120, 144, 168, 192, 216, 240, 264, 288, 312, 336, 360, 384, 408, 432, 456, 480, 504, 528, 552, 576, 600, 624, 648, 672, 696, 720, 744, 768, 792, 816, 840, 864, 888, 912, 936, 960, 984, 1008, 1032, 1056, 1080, 1104, 1128, 1152, 1176, 1200, 1224, 1248, 1272, 1296, 1320, 1344, 1368, 1392, 1416, 1440, 1464, 1488, 1512, 1536, 1560, 1584, 1608, 1632, 1656, 1680, 1704, 1728, 1752, 1776, 1800, 1824, 1848, 1872, 1896, 1920, 1944, 1968, 1992, 2016, 2040, 2064, 2088, 2112, 2136, 2160, 2184, 2208, 2232, 2256, 2280, 2304, 2328, 2352, 2376, 2400, 2424, 2448, 2472, 2496, 2520, 2544, 2568, 2592, 2616, 2640, 2664, 2688, 2712, 2736, 2760, 2784, 2808, 2832, 2856, 2880, 2904, 2928, 2952, 2976, 3000, 3024, 3048, 3072, 3096, 3120, 3144, 3168, 3192, 3216, 3240, 3264, 3288, 3312, 3336, 3360, 3384, 3408, 3432, 3456, 3480, 3504, 3528, 3552, 3576, 3600, 3624, 3648, 3672, 3696, 3720, 3744, 3768, 3792, 3816, 3840, 3864, 3888, 3912, 3936, 3960, 3984, 4008, 4032, 4056, 4080, 4104, 4128, 4152, 4176, 4200, 4224, 4248, 4272, 4296, 4320, 4344, 4368, 4392, 4416, 4440, 4464, 4488, 4512, 4536, 4560, 4584, 4608, 4632, 4656, 4680, 4704, 4728, 4752, 4776, 4800, 4824, 4848, 4872, 4896, 4920, 4944, 4968, 4992, 5016, 5040, 5064, 5088, 5112, 5136, 5160, 5184, 5208, 5232, 5256, 5280, 5304, 5328, 5352, 5376, 5400, 5424, 5448, 5472, 5496, 5520, 5544, 5568, 5592, 5616, 5640, 5664, 5688, 5712, 5736, 5760, 5784, 5808, 5832, 5856, 5880, 5904, 5928, 5952, 5976, 6000, 6024, 6048, 6072, 6096, 6120, 
0, 25, 50, 75, 100, 125, 150, 175, 200, 225, 250, 275, 300, 325, 350, 375, 400, 425, 450, 475, 500, 525, 550, 575, 600, 625, 650, 675, 700, 725, 750, 775, 800, 825, 850, 875, 900, 925, 950, 975, 1000, 1025, 1050, 1075, 1100, 1125, 1150, 1175, 1200, 1225, 1250, 1275, 1300, 1325, 1350, 1375, 1400, 1425, 1450, 1475, 1500, 1525, 1550, 1575, 1600, 1625, 1650, 1675, 1700, 1725, 1750, 1775, 1800, 1825, 1850, 1875, 1900, 1925, 1950, 1975, 2000, 2025, 2050, 2075, 2100, 2125, 2150, 2175, 2200, 2225, 2250, 2275, 2300, 2325, 2350, 2375, 2400, 2425, 2450, 2475, 2500, 2525, 2550, 2575, 2600, 2625, 2650, 2675, 2700, 2725, 2750, 2775, 2800, 2825, 2850, 2875, 2900, 2925, 2950, 2975, 3000, 3025, 3050, 3075, 3100, 3125, 3150, 3175, 3200, 3225, 3250, 3275, 3300, 3325, 3350, 3375, 3400, 3425, 3450, 3475, 3500, 3525, 3550, 3575, 3600, 3625, 3650, 3675, 3700, 3725, 3750, 3775, 3800, 3825, 3850, 3875, 3900, 3925, 3950, 3975, 4000, 4025, 4050, 4075, 4100, 4125, 4150, 4175, 4200, 4225, 4250, 4275, 4300, 4325, 4350, 4375, 4400, 4425, 4450, 4475, 4500, 4525, 4550, 4575, 4600, 4625, 4650, 4675, 4700, 4725, 4750, 4775, 4800, 4825, 4850, 4875, 4900, 4925, 4950, 4975, 5000, 5025, 5050, 5075, 5100, 5125, 5150, 5175, 5200, 5225, 5250, 5275, 5300, 5325, 5350, 5375, 5400, 5425, 5450, 5475, 5500, 5525, 5550, 5575, 5600, 5625, 5650, 5675, 5700, 5725, 5750, 5775, 5800, 5825, 5850, 5875, 5900, 5925, 5950, 5975, 6000, 6025, 6050, 6075, 6100, 6125, 6150, 6175, 6200, 6225, 6250, 6275, 6300, 6325, 6350, 6375, 
0, 26, 52, 78, 104, 130, 156, 182, 208, 234, 260, 286, 312, 338, 364, 390, 416, 442, 468, 494, 520, 546, 572, 598, 624, 650, 676, 702, 728, 754, 780, 806, 832, 858, 884, 910, 936, 962, 988, 1014, 1040, 1066, 1092, 1118, 1144, 1170, 1196, 1222, 1248, 1274, 1300, 1326, 1352, 1378, 1404, 1430, 1456, 1482, 1508, 1534, 1560, 1586, 1612, 1638, 1664, 1690, 1716, 1742, 1768, 1794, 1820, 1846, 1872, 1898, 1924, 1950, 1976, 2002, 2028, 2054, 2080, 2106, 2132, 2158, 2184, 2210, 2236, 2262, 2288, 2314, 2340, 2366, 2392, 2418, 2444, 2470, 2496, 2522, 2548, 2574, 2600, 2626, 2652, 2678, 2704, 2730, 2756, 2782, 2808, 2834, 2860, 2886, 2912, 2938, 2964, 2990, 3016, 3042, 3068, 3094, 3120, 3146, 3172, 3198, 3224, 3250, 3276, 3302, 3328, 3354, 3380, 3406, 3432, 3458, 3484, 3510, 3536, 3562, 3588, 3614, 3640, 3666, 3692, 3718, 3744, 3770, 3796, 3822, 3848, 3874, 3900, 3926, 3952, 3978, 4004, 4030, 4056, 4082, 4108, 4134, 4160, 4186, 4212, 4238, 4264, 4290, 4316, 4342, 4368, 4394, 4420, 4446, 4472, 4498, 4524, 4550, 4576, 4602, 4628, 4654, 4680, 4706, 4732, 4758, 4784, 4810, 4836, 4862, 4888, 4914, 4940, 4966, 4992, 5018, 5044, 5070, 5096, 5122, 5148, 5174, 5200, 5226, 5252, 5278, 5304, 5330, 5356, 5382, 5408, 5434, 5460, 5486, 5512, 5538, 5564, 5590, 5616, 5642, 5668, 5694, 5720, 5746, 5772, 5798, 5824, 5850, 5876, 5902, 5928, 5954, 5980, 6006, 6032, 6058, 6084, 6110, 6136, 6162, 6188, 6214, 6240, 6266, 6292, 6318, 6344, 6370, 6396, 6422, 6448, 6474, 6500, 6526, 6552, 6578, 6604, 6630, 
0, 27, 54, 81, 108, 135, 162, 189, 216, 243, 270, 297, 324, 351, 378, 405, 432, 459, 486, 513, 540, 567, 594, 621, 648, 675, 702, 729, 756, 783, 810, 837, 864, 891, 918, 945, 972, 999, 1026, 1053, 1080, 1107, 1134, 1161, 1188, 1215, 1242, 1269, 1296, 1323, 1350, 1377, 1404, 1431, 1458, 1485, 1512, 1539, 1566, 1593, 1620, 1647, 1674, 1701, 1728, 1755, 1782, 1809, 1836, 1863, 1890, 1917, 1944, 1971, 1998, 2025, 2052, 2079, 2106, 2133, 2160, 2187, 2214, 2241, 2268, 2295, 2322, 2349, 2376, 2403, 2430, 2457, 2484, 2511, 2538, 2565, 2592, 2619, 2646, 2673, 2700, 2727, 2754, 2781, 2808, 2835, 2862, 2889, 2916, 2943, 2970, 2997, 3024, 3051, 3078, 3105, 3132, 3159, 3186, 3213, 3240, 3267, 3294, 3321, 3348, 3375, 3402, 3429, 3456, 3483, 3510, 3537, 3564, 3591, 3618, 3645, 3672, 3699, 3726, 3753, 3780, 3807, 3834, 3861, 3888, 3915, 3942, 3969, 3996, 4023, 4050, 4077, 4104, 4131, 4158, 4185, 4212, 4239, 4266, 4293, 4320, 4347, 4374, 4401, 4428, 4455, 4482, 4509, 4536, 4563, 4590, 4617, 4644, 4671, 4698, 4725, 4752, 4779, 4806, 4833, 4860, 4887, 4914, 4941, 4968, 4995, 5022, 5049, 5076, 5103, 5130, 5157, 5184, 5211, 5238, 5265, 5292, 5319, 5346, 5373, 5400, 5427, 5454, 5481, 5508, 5535, 5562, 5589, 5616, 5643, 5670, 5697, 5724, 5751, 5778, 5805, 5832, 5859, 5886, 5913, 5940, 5967, 5994, 6021, 6048, 6075, 6102, 6129, 6156, 6183, 6210, 6237, 6264, 6291, 6318, 6345, 6372, 6399, 6426, 6453, 6480, 6507, 6534, 6561, 6588, 6615, 6642, 6669, 6696, 6723, 6750, 6777, 6804, 6831, 6858, 6885, 
0, 28, 56, 84, 112, 140, 168, 196, 224, 252, 280, 308, 336, 364, 392, 420, 448, 476, 504, 532, 560, 588, 616, 644, 672, 700, 728, 756, 784, 812, 840, 868, 896, 924, 952, 980, 1008, 1036, 1064, 1092, 1120, 1148, 1176, 1204, 1232, 1260, 1288, 1316, 1344, 1372, 1400, 1428, 1456, 1484, 1512, 1540, 1568, 1596, 1624, 1652, 1680, 1708, 1736, 1764, 1792, 1820, 1848, 1876, 1904, 1932, 1960, 1988, 2016, 2044, 2072, 2100, 2128, 2156, 2184, 2212, 2240, 2268, 2296, 2324, 2352, 2380, 2408, 2436, 2464, 2492, 2520, 2548, 2576, 2604, 2632, 2660, 2688, 2716, 2744, 2772, 2800, 2828, 2856, 2884, 2912, 2940, 2968, 2996, 3024, 3052, 3080, 3108, 3136, 3164, 3192, 3220, 3248, 3276, 3304, 3332, 3360, 3388, 3416, 3444, 3472, 3500, 3528, 3556, 3584, 3612, 3640, 3668, 3696, 3724, 3752, 3780, 3808, 3836, 3864, 3892, 3920, 3948, 3976, 4004, 4032, 4060, 4088, 4116, 4144, 4172, 4200, 4228, 4256, 4284, 4312, 4340, 4368, 4396, 4424, 4452, 4480, 4508, 4536, 4564, 4592, 4620, 4648, 4676, 4704, 4732, 4760, 4788, 4816, 4844, 4872, 4900, 4928, 4956, 4984, 5012, 5040, 5068, 5096, 5124, 5152, 5180, 5208, 5236, 5264, 5292, 5320, 5348, 5376, 5404, 5432, 5460, 5488, 5516, 5544, 5572, 5600, 5628, 5656, 5684, 5712, 5740, 5768, 5796, 5824, 5852, 5880, 5908, 5936, 5964, 5992, 6020, 6048, 6076, 6104, 6132, 6160, 6188, 6216, 6244, 6272, 6300, 6328, 6356, 6384, 6412, 6440, 6468, 6496, 6524, 6552, 6580, 6608, 6636, 6664, 6692, 6720, 6748, 6776, 6804, 6832, 6860, 6888, 6916, 6944, 6972, 7000, 7028, 7056, 7084, 7112, 7140, 
0, 29, 58, 87, 116, 145, 174, 203, 232, 261, 290, 319, 348, 377, 406, 435, 464, 493, 522, 551, 580, 609, 638, 667, 696, 725, 754, 783, 812, 841, 870, 899, 928, 957, 986, 1015, 1044, 1073, 1102, 1131, 1160, 1189, 1218, 1247, 1276, 1305, 1334, 1363, 1392, 1421, 1450, 1479, 1508, 1537, 1566, 1595, 1624, 1653, 1682, 1711, 1740, 1769, 1798, 1827, 1856, 1885, 1914, 1943, 1972, 2001, 2030, 2059, 2088, 2117, 2146, 2175, 2204, 2233, 2262, 2291, 2320, 2349, 2378, 2407, 2436, 2465, 2494, 2523, 2552, 2581, 2610, 2639, 2668, 2697, 2726, 2755, 2784, 2813, 2842, 2871, 2900, 2929, 2958, 2987, 3016, 3045, 3074, 3103, 3132, 3161, 3190, 3219, 3248, 3277, 3306, 3335, 3364, 3393, 3422, 3451, 3480, 3509, 3538, 3567, 3596, 3625, 3654, 3683, 3712, 3741, 3770, 3799, 3828, 3857, 3886, 3915, 3944, 3973, 4002, 4031, 4060, 4089, 4118, 4147, 4176, 4205, 4234, 4263, 4292, 4321, 4350, 4379, 4408, 4437, 4466, 4495, 4524, 4553, 4582, 4611, 4640, 4669, 4698, 4727, 4756, 4785, 4814, 4843, 4872, 4901, 4930, 4959, 4988, 5017, 5046, 5075, 5104, 5133, 5162, 5191, 5220, 5249, 5278, 5307, 5336, 5365, 5394, 5423, 5452, 5481, 5510, 5539, 5568, 5597, 5626, 5655, 5684, 5713, 5742, 5771, 5800, 5829, 5858, 5887, 5916, 5945, 5974, 6003, 6032, 6061, 6090, 6119, 6148, 6177, 6206, 6235, 6264, 6293, 6322, 6351, 6380, 6409, 6438, 6467, 6496, 6525, 6554, 6583, 6612, 6641, 6670, 6699, 6728, 6757, 6786, 6815, 6844, 6873, 6902, 6931, 6960, 6989, 7018, 7047, 7076, 7105, 7134, 7163, 7192, 7221, 7250, 7279, 7308, 7337, 7366, 7395, 
0, 30, 60, 90, 120, 150, 180, 210, 240, 270, 300, 330, 360, 390, 420, 450, 480, 510, 540, 570, 600, 630, 660, 690, 720, 750, 780, 810, 840, 870, 900, 930, 960, 990, 1020, 1050, 1080, 1110, 1140, 1170, 1200, 1230, 1260, 1290, 1320, 1350, 1380, 1410, 1440, 1470, 1500, 1530, 1560, 1590, 1620, 1650, 1680, 1710, 1740, 1770, 1800, 1830, 1860, 1890, 1920, 1950, 1980, 2010, 2040, 2070, 2100, 2130, 2160, 2190, 2220, 2250, 2280, 2310, 2340, 2370, 2400, 2430, 2460, 2490, 2520, 2550, 2580, 2610, 2640, 2670, 2700, 2730, 2760, 2790, 2820, 2850, 2880, 2910, 2940, 2970, 3000, 3030, 3060, 3090, 3120, 3150, 3180, 3210, 3240, 3270, 3300, 3330, 3360, 3390, 3420, 3450, 3480, 3510, 3540, 3570, 3600, 3630, 3660, 3690, 3720, 3750, 3780, 3810, 3840, 3870, 3900, 3930, 3960, 3990, 4020, 4050, 4080, 4110, 4140, 4170, 4200, 4230, 4260, 4290, 4320, 4350, 4380, 4410, 4440, 4470, 4500, 4530, 4560, 4590, 4620, 4650, 4680, 4710, 4740, 4770, 4800, 4830, 4860, 4890, 4920, 4950, 4980, 5010, 5040, 5070, 5100, 5130, 5160, 5190, 5220, 5250, 5280, 5310, 5340, 5370, 5400, 5430, 5460, 5490, 5520, 5550, 5580, 5610, 5640, 5670, 5700, 5730, 5760, 5790, 5820, 5850, 5880, 5910, 5940, 5970, 6000, 6030, 6060, 6090, 6120, 6150, 6180, 6210, 6240, 6270, 6300, 6330, 6360, 6390, 6420, 6450, 6480, 6510, 6540, 6570, 6600, 6630, 6660, 6690, 6720, 6750, 6780, 6810, 6840, 6870, 6900, 6930, 6960, 6990, 7020, 7050, 7080, 7110, 7140, 7170, 7200, 7230, 7260, 7290, 7320, 7350, 7380, 7410, 7440, 7470, 7500, 7530, 7560, 7590, 7620, 7650, 
0, 31, 62, 93, 124, 155, 186, 217, 248, 279, 310, 341, 372, 403, 434, 465, 496, 527, 558, 589, 620, 651, 682, 713, 744, 775, 806, 837, 868, 899, 930, 961, 992, 1023, 1054, 1085, 1116, 1147, 1178, 1209, 1240, 1271, 1302, 1333, 1364, 1395, 1426, 1457, 1488, 1519, 1550, 1581, 1612, 1643, 1674, 1705, 1736, 1767, 1798, 1829, 1860, 1891, 1922, 1953, 1984, 2015, 2046, 2077, 2108, 2139, 2170, 2201, 2232, 2263, 2294, 2325, 2356, 2387, 2418, 2449, 2480, 2511, 2542, 2573, 2604, 2635, 2666, 2697, 2728, 2759, 2790, 2821, 2852, 2883, 2914, 2945, 2976, 3007, 3038, 3069, 3100, 3131, 3162, 3193, 3224, 3255, 3286, 3317, 3348, 3379, 3410, 3441, 3472, 3503, 3534, 3565, 3596, 3627, 3658, 3689, 3720, 3751, 3782, 3813, 3844, 3875, 3906, 3937, 3968, 3999, 4030, 4061, 4092, 4123, 4154, 4185, 4216, 4247, 4278, 4309, 4340, 4371, 4402, 4433, 4464, 4495, 4526, 4557, 4588, 4619, 4650, 4681, 4712, 4743, 4774, 4805, 4836, 4867, 4898, 4929, 4960, 4991, 5022, 5053, 5084, 5115, 5146, 5177, 5208, 5239, 5270, 5301, 5332, 5363, 5394, 5425, 5456, 5487, 5518, 5549, 5580, 5611, 5642, 5673, 5704, 5735, 5766, 5797, 5828, 5859, 5890, 5921, 5952, 5983, 6014, 6045, 6076, 6107, 6138, 6169, 6200, 6231, 6262, 6293, 6324, 6355, 6386, 6417, 6448, 6479, 6510, 6541, 6572, 6603, 6634, 6665, 6696, 6727, 6758, 6789, 6820, 6851, 6882, 6913, 6944, 6975, 7006, 7037, 7068, 7099, 7130, 7161, 7192, 7223, 7254, 7285, 7316, 7347, 7378, 7409, 7440, 7471, 7502, 7533, 7564, 7595, 7626, 7657, 7688, 7719, 7750, 7781, 7812, 7843, 7874, 7905, 
0, 32, 64, 96, 128, 160, 192, 224, 256, 288, 320, 352, 384, 416, 448, 480, 512, 544, 576, 608, 640, 672, 704, 736, 768, 800, 832, 864, 896, 928, 960, 992, 1024, 1056, 1088, 1120, 1152, 1184, 1216, 1248, 1280, 1312, 1344, 1376, 1408, 1440, 1472, 1504, 1536, 1568, 1600, 1632, 1664, 1696, 1728, 1760, 1792, 1824, 1856, 1888, 1920, 1952, 1984, 2016, 2048, 2080, 2112, 2144, 2176, 2208, 2240, 2272, 2304, 2336, 2368, 2400, 2432, 2464, 2496, 2528, 2560, 2592, 2624, 2656, 2688, 2720, 2752, 2784, 2816, 2848, 2880, 2912, 2944, 2976, 3008, 3040, 3072, 3104, 3136, 3168, 3200, 3232, 3264, 3296, 3328, 3360, 3392, 3424, 3456, 3488, 3520, 3552, 3584, 3616, 3648, 3680, 3712, 3744, 3776, 3808, 3840, 3872, 3904, 3936, 3968, 4000, 4032, 4064, 4096, 4128, 4160, 4192, 4224, 4256, 4288, 4320, 4352, 4384, 4416, 4448, 4480, 4512, 4544, 4576, 4608, 4640, 4672, 4704, 4736, 4768, 4800, 4832, 4864, 4896, 4928, 4960, 4992, 5024, 5056, 5088, 5120, 5152, 5184, 5216, 5248, 5280, 5312, 5344, 5376, 5408, 5440, 5472, 5504, 5536, 5568, 5600, 5632, 5664, 5696, 5728, 5760, 5792, 5824, 5856, 5888, 5920, 5952, 5984, 6016, 6048, 6080, 6112, 6144, 6176, 6208, 6240, 6272, 6304, 6336, 6368, 6400, 6432, 6464, 6496, 6528, 6560, 6592, 6624, 6656, 6688, 6720, 6752, 6784, 6816, 6848, 6880, 6912, 6944, 6976, 7008, 7040, 7072, 7104, 7136, 7168, 7200, 7232, 7264, 7296, 7328, 7360, 7392, 7424, 7456, 7488, 7520, 7552, 7584, 7616, 7648, 7680, 7712, 7744, 7776, 7808, 7840, 7872, 7904, 7936, 7968, 8000, 8032, 8064, 8096, 8128, 8160, 
0, 33, 66, 99, 132, 165, 198, 231, 264, 297, 330, 363, 396, 429, 462, 495, 528, 561, 594, 627, 660, 693, 726, 759, 792, 825, 858, 891, 924, 957, 990, 1023, 1056, 1089, 1122, 1155, 1188, 1221, 1254, 1287, 1320, 1353, 1386, 1419, 1452, 1485, 1518, 1551, 1584, 1617, 1650, 1683, 1716, 1749, 1782, 1815, 1848, 1881, 1914, 1947, 1980, 2013, 2046, 2079, 2112, 2145, 2178, 2211, 2244, 2277, 2310, 2343, 2376, 2409, 2442, 2475, 2508, 2541, 2574, 2607, 2640, 2673, 2706, 2739, 2772, 2805, 2838, 2871, 2904, 2937, 2970, 3003, 3036, 3069, 3102, 3135, 3168, 3201, 3234, 3267, 3300, 3333, 3366, 3399, 3432, 3465, 3498, 3531, 3564, 3597, 3630, 3663, 3696, 3729, 3762, 3795, 3828, 3861, 3894, 3927, 3960, 3993, 4026, 4059, 4092, 4125, 4158, 4191, 4224, 4257, 4290, 4323, 4356, 4389, 4422, 4455, 4488, 4521, 4554, 4587, 4620, 4653, 4686, 4719, 4752, 4785, 4818, 4851, 4884, 4917, 4950, 4983, 5016, 5049, 5082, 5115, 5148, 5181, 5214, 5247, 5280, 5313, 5346, 5379, 5412, 5445, 5478, 5511, 5544, 5577, 5610, 5643, 5676, 5709, 5742, 5775, 5808, 5841, 5874, 5907, 5940, 5973, 6006, 6039, 6072, 6105, 6138, 6171, 6204, 6237, 6270, 6303, 6336, 6369, 6402, 6435, 6468, 6501, 6534, 6567, 6600, 6633, 6666, 6699, 6732, 6765, 6798, 6831, 6864, 6897, 6930, 6963, 6996, 7029, 7062, 7095, 7128, 7161, 7194, 7227, 7260, 7293, 7326, 7359, 7392, 7425, 7458, 7491, 7524, 7557, 7590, 7623, 7656, 7689, 7722, 7755, 7788, 7821, 7854, 7887, 7920, 7953, 7986, 8019, 8052, 8085, 8118, 8151, 8184, 8217, 8250, 8283, 8316, 8349, 8382, 8415, 
0, 34, 68, 102, 136, 170, 204, 238, 272, 306, 340, 374, 408, 442, 476, 510, 544, 578, 612, 646, 680, 714, 748, 782, 816, 850, 884, 918, 952, 986, 1020, 1054, 1088, 1122, 1156, 1190, 1224, 1258, 1292, 1326, 1360, 1394, 1428, 1462, 1496, 1530, 1564, 1598, 1632, 1666, 1700, 1734, 1768, 1802, 1836, 1870, 1904, 1938, 1972, 2006, 2040, 2074, 2108, 2142, 2176, 2210, 2244, 2278, 2312, 2346, 2380, 2414, 2448, 2482, 2516, 2550, 2584, 2618, 2652, 2686, 2720, 2754, 2788, 2822, 2856, 2890, 2924, 2958, 2992, 3026, 3060, 3094, 3128, 3162, 3196, 3230, 3264, 3298, 3332, 3366, 3400, 3434, 3468, 3502, 3536, 3570, 3604, 3638, 3672, 3706, 3740, 3774, 3808, 3842, 3876, 3910, 3944, 3978, 4012, 4046, 4080, 4114, 4148, 4182, 4216, 4250, 4284, 4318, 4352, 4386, 4420, 4454, 4488, 4522, 4556, 4590, 4624, 4658, 4692, 4726, 4760, 4794, 4828, 4862, 4896, 4930, 4964, 4998, 5032, 5066, 5100, 5134, 5168, 5202, 5236, 5270, 5304, 5338, 5372, 5406, 5440, 5474, 5508, 5542, 5576, 5610, 5644, 5678, 5712, 5746, 5780, 5814, 5848, 5882, 5916, 5950, 5984, 6018, 6052, 6086, 6120, 6154, 6188, 6222, 6256, 6290, 6324, 6358, 6392, 6426, 6460, 6494, 6528, 6562, 6596, 6630, 6664, 6698, 6732, 6766, 6800, 6834, 6868, 6902, 6936, 6970, 7004, 7038, 7072, 7106, 7140, 7174, 7208, 7242, 7276, 7310, 7344, 7378, 7412, 7446, 7480, 7514, 7548, 7582, 7616, 7650, 7684, 7718, 7752, 7786, 7820, 7854, 7888, 7922, 7956, 7990, 8024, 8058, 8092, 8126, 8160, 8194, 8228, 8262, 8296, 8330, 8364, 8398, 8432, 8466, 8500, 8534, 8568, 8602, 8636, 8670, 
0, 35, 70, 105, 140, 175, 210, 245, 280, 315, 350, 385, 420, 455, 490, 525, 560, 595, 630, 665, 700, 735, 770, 805, 840, 875, 910, 945, 980, 1015, 1050, 1085, 1120, 1155, 1190, 1225, 1260, 1295, 1330, 1365, 1400, 1435, 1470, 1505, 1540, 1575, 1610, 1645, 1680, 1715, 1750, 1785, 1820, 1855, 1890, 1925, 1960, 1995, 2030, 2065, 2100, 2135, 2170, 2205, 2240, 2275, 2310, 2345, 2380, 2415, 2450, 2485, 2520, 2555, 2590, 2625, 2660, 2695, 2730, 2765, 2800, 2835, 2870, 2905, 2940, 2975, 3010, 3045, 3080, 3115, 3150, 3185, 3220, 3255, 3290, 3325, 3360, 3395, 3430, 3465, 3500, 3535, 3570, 3605, 3640, 3675, 3710, 3745, 3780, 3815, 3850, 3885, 3920, 3955, 3990, 4025, 4060, 4095, 4130, 4165, 4200, 4235, 4270, 4305, 4340, 4375, 4410, 4445, 4480, 4515, 4550, 4585, 4620, 4655, 4690, 4725, 4760, 4795, 4830, 4865, 4900, 4935, 4970, 5005, 5040, 5075, 5110, 5145, 5180, 5215, 5250, 5285, 5320, 5355, 5390, 5425, 5460, 5495, 5530, 5565, 5600, 5635, 5670, 5705, 5740, 5775, 5810, 5845, 5880, 5915, 5950, 5985, 6020, 6055, 6090, 6125, 6160, 6195, 6230, 6265, 6300, 6335, 6370, 6405, 6440, 6475, 6510, 6545, 6580, 6615, 6650, 6685, 6720, 6755, 6790, 6825, 6860, 6895, 6930, 6965, 7000, 7035, 7070, 7105, 7140, 7175, 7210, 7245, 7280, 7315, 7350, 7385, 7420, 7455, 7490, 7525, 7560, 7595, 7630, 7665, 7700, 7735, 7770, 7805, 7840, 7875, 7910, 7945, 7980, 8015, 8050, 8085, 8120, 8155, 8190, 8225, 8260, 8295, 8330, 8365, 8400, 8435, 8470, 8505, 8540, 8575, 8610, 8645, 8680, 8715, 8750, 8785, 8820, 8855, 8890, 8925, 
0, 36, 72, 108, 144, 180, 216, 252, 288, 324, 360, 396, 432, 468, 504, 540, 576, 612, 648, 684, 720, 756, 792, 828, 864, 900, 936, 972, 1008, 1044, 1080, 1116, 1152, 1188, 1224, 1260, 1296, 1332, 1368, 1404, 1440, 1476, 1512, 1548, 1584, 1620, 1656, 1692, 1728, 1764, 1800, 1836, 1872, 1908, 1944, 1980, 2016, 2052, 2088, 2124, 2160, 2196, 2232, 2268, 2304, 2340, 2376, 2412, 2448, 2484, 2520, 2556, 2592, 2628, 2664, 2700, 2736, 2772, 2808, 2844, 2880, 2916, 2952, 2988, 3024, 3060, 3096, 3132, 3168, 3204, 3240, 3276, 3312, 3348, 3384, 3420, 3456, 3492, 3528, 3564, 3600, 3636, 3672, 3708, 3744, 3780, 3816, 3852, 3888, 3924, 3960, 3996, 4032, 4068, 4104, 4140, 4176, 4212, 4248, 4284, 4320, 4356, 4392, 4428, 4464, 4500, 4536, 4572, 4608, 4644, 4680, 4716, 4752, 4788, 4824, 4860, 4896, 4932, 4968, 5004, 5040, 5076, 5112, 5148, 5184, 5220, 5256, 5292, 5328, 5364, 5400, 5436, 5472, 5508, 5544, 5580, 5616, 5652, 5688, 5724, 5760, 5796, 5832, 5868, 5904, 5940, 5976, 6012, 6048, 6084, 6120, 6156, 6192, 6228, 6264, 6300, 6336, 6372, 6408, 6444, 6480, 6516, 6552, 6588, 6624, 6660, 6696, 6732, 6768, 6804, 6840, 6876, 6912, 6948, 6984, 7020, 7056, 7092, 7128, 7164, 7200, 7236, 7272, 7308, 7344, 7380, 7416, 7452, 7488, 7524, 7560, 7596, 7632, 7668, 7704, 7740, 7776, 7812, 7848, 7884, 7920, 7956, 7992, 8028, 8064, 8100, 8136, 8172, 8208, 8244, 8280, 8316, 8352, 8388, 8424, 8460, 8496, 8532, 8568, 8604, 8640, 8676, 8712, 8748, 8784, 8820, 8856, 8892, 8928, 8964, 9000, 9036, 9072, 9108, 9144, 9180, 
0, 37, 74, 111, 148, 185, 222, 259, 296, 333, 370, 407, 444, 481, 518, 555, 592, 629, 666, 703, 740, 777, 814, 851, 888, 925, 962, 999, 1036, 1073, 1110, 1147, 1184, 1221, 1258, 1295, 1332, 1369, 1406, 1443, 1480, 1517, 1554, 1591, 1628, 1665, 1702, 1739, 1776, 1813, 1850, 1887, 1924, 1961, 1998, 2035, 2072, 2109, 2146, 2183, 2220, 2257, 2294, 2331, 2368, 2405, 2442, 2479, 2516, 2553, 2590, 2627, 2664, 2701, 2738, 2775, 2812, 2849, 2886, 2923, 2960, 2997, 3034, 3071, 3108, 3145, 3182, 3219, 3256, 3293, 3330, 3367, 3404, 3441, 3478, 3515, 3552, 3589, 3626, 3663, 3700, 3737, 3774, 3811, 3848, 3885, 3922, 3959, 3996, 4033, 4070, 4107, 4144, 4181, 4218, 4255, 4292, 4329, 4366, 4403, 4440, 4477, 4514, 4551, 4588, 4625, 4662, 4699, 4736, 4773, 4810, 4847, 4884, 4921, 4958, 4995, 5032, 5069, 5106, 5143, 5180, 5217, 5254, 5291, 5328, 5365, 5402, 5439, 5476, 5513, 5550, 5587, 5624, 5661, 5698, 5735, 5772, 5809, 5846, 5883, 5920, 5957, 5994, 6031, 6068, 6105, 6142, 6179, 6216, 6253, 6290, 6327, 6364, 6401, 6438, 6475, 6512, 6549, 6586, 6623, 6660, 6697, 6734, 6771, 6808, 6845, 6882, 6919, 6956, 6993, 7030, 7067, 7104, 7141, 7178, 7215, 7252, 7289, 7326, 7363, 7400, 7437, 7474, 7511, 7548, 7585, 7622, 7659, 7696, 7733, 7770, 7807, 7844, 7881, 7918, 7955, 7992, 8029, 8066, 8103, 8140, 8177, 8214, 8251, 8288, 8325, 8362, 8399, 8436, 8473, 8510, 8547, 8584, 8621, 8658, 8695, 8732, 8769, 8806, 8843, 8880, 8917, 8954, 8991, 9028, 9065, 9102, 9139, 9176, 9213, 9250, 9287, 9324, 9361, 9398, 9435, 
0, 38, 76, 114, 152, 190, 228, 266, 304, 342, 380, 418, 456, 494, 532, 570, 608, 646, 684, 722, 760, 798, 836, 874, 912, 950, 988, 1026, 1064, 1102, 1140, 1178, 1216, 1254, 1292, 1330, 1368, 1406, 1444, 1482, 1520, 1558, 1596, 1634, 1672, 1710, 1748, 1786, 1824, 1862, 1900, 1938, 1976, 2014, 2052, 2090, 2128, 2166, 2204, 2242, 2280, 2318, 2356, 2394, 2432, 2470, 2508, 2546, 2584, 2622, 2660, 2698, 2736, 2774, 2812, 2850, 2888, 2926, 2964, 3002, 3040, 3078, 3116, 3154, 3192, 3230, 3268, 3306, 3344, 3382, 3420, 3458, 3496, 3534, 3572, 3610, 3648, 3686, 3724, 3762, 3800, 3838, 3876, 3914, 3952, 3990, 4028, 4066, 4104, 4142, 4180, 4218, 4256, 4294, 4332, 4370, 4408, 4446, 4484, 4522, 4560, 4598, 4636, 4674, 4712, 4750, 4788, 4826, 4864, 4902, 4940, 4978, 5016, 5054, 5092, 5130, 5168, 5206, 5244, 5282, 5320, 5358, 5396, 5434, 5472, 5510, 5548, 5586, 5624, 5662, 5700, 5738, 5776, 5814, 5852, 5890, 5928, 5966, 6004, 6042, 6080, 6118, 6156, 6194, 6232, 6270, 6308, 6346, 6384, 6422, 6460, 6498, 6536, 6574, 6612, 6650, 6688, 6726, 6764, 6802, 6840, 6878, 6916, 6954, 6992, 7030, 7068, 7106, 7144, 7182, 7220, 7258, 7296, 7334, 7372, 7410, 7448, 7486, 7524, 7562, 7600, 7638, 7676, 7714, 7752, 7790, 7828, 7866, 7904, 7942, 7980, 8018, 8056, 8094, 8132, 8170, 8208, 8246, 8284, 8322, 8360, 8398, 8436, 8474, 8512, 8550, 8588, 8626, 8664, 8702, 8740, 8778, 8816, 8854, 8892, 8930, 8968, 9006, 9044, 9082, 9120, 9158, 9196, 9234, 9272, 9310, 9348, 9386, 9424, 9462, 9500, 9538, 9576, 9614, 9652, 9690, 
0, 39, 78, 117, 156, 195, 234, 273, 312, 351, 390, 429, 468, 507, 546, 585, 624, 663, 702, 741, 780, 819, 858, 897, 936, 975, 1014, 1053, 1092, 1131, 1170, 1209, 1248, 1287, 1326, 1365, 1404, 1443, 1482, 1521, 1560, 1599, 1638, 1677, 1716, 1755, 1794, 1833, 1872, 1911, 1950, 1989, 2028, 2067, 2106, 2145, 2184, 2223, 2262, 2301, 2340, 2379, 2418, 2457, 2496, 2535, 2574, 2613, 2652, 2691, 2730, 2769, 2808, 2847, 2886, 2925, 2964, 3003, 3042, 3081, 3120, 3159, 3198, 3237, 3276, 3315, 3354, 3393, 3432, 3471, 3510, 3549, 3588, 3627, 3666, 3705, 3744, 3783, 3822, 3861, 3900, 3939, 3978, 4017, 4056, 4095, 4134, 4173, 4212, 4251, 4290, 4329, 4368, 4407, 4446, 4485, 4524, 4563, 4602, 4641, 4680, 4719, 4758, 4797, 4836, 4875, 4914, 4953, 4992, 5031, 5070, 5109, 5148, 5187, 5226, 5265, 5304, 5343, 5382, 5421, 5460, 5499, 5538, 5577, 5616, 5655, 5694, 5733, 5772, 5811, 5850, 5889, 5928, 5967, 6006, 6045, 6084, 6123, 6162, 6201, 6240, 6279, 6318, 6357, 6396, 6435, 6474, 6513, 6552, 6591, 6630, 6669, 6708, 6747, 6786, 6825, 6864, 6903, 6942, 6981, 7020, 7059, 7098, 7137, 7176, 7215, 7254, 7293, 7332, 7371, 7410, 7449, 7488, 7527, 7566, 7605, 7644, 7683, 7722, 7761, 7800, 7839, 7878, 7917, 7956, 7995, 8034, 8073, 8112, 8151, 8190, 8229, 8268, 8307, 8346, 8385, 8424, 8463, 8502, 8541, 8580, 8619, 8658, 8697, 8736, 8775, 8814, 8853, 8892, 8931, 8970, 9009, 9048, 9087, 9126, 9165, 9204, 9243, 9282, 9321, 9360, 9399, 9438, 9477, 9516, 9555, 9594, 9633, 9672, 9711, 9750, 9789, 9828, 9867, 9906, 9945, 
0, 40, 80, 120, 160, 200, 240, 280, 320, 360, 400, 440, 480, 520, 560, 600, 640, 680, 720, 760, 800, 840, 880, 920, 960, 1000, 1040, 1080, 1120, 1160, 1200, 1240, 1280, 1320, 1360, 1400, 1440, 1480, 1520, 1560, 1600, 1640, 1680, 1720, 1760, 1800, 1840, 1880, 1920, 1960, 2000, 2040, 2080, 2120, 2160, 2200, 2240, 2280, 2320, 2360, 2400, 2440, 2480, 2520, 2560, 2600, 2640, 2680, 2720, 2760, 2800, 2840, 2880, 2920, 2960, 3000, 3040, 3080, 3120, 3160, 3200, 3240, 3280, 3320, 3360, 3400, 3440, 3480, 3520, 3560, 3600, 3640, 3680, 3720, 3760, 3800, 3840, 3880, 3920, 3960, 4000, 4040, 4080, 4120, 4160, 4200, 4240, 4280, 4320, 4360, 4400, 4440, 4480, 4520, 4560, 4600, 4640, 4680, 4720, 4760, 4800, 4840, 4880, 4920, 4960, 5000, 5040, 5080, 5120, 5160, 5200, 5240, 5280, 5320, 5360, 5400, 5440, 5480, 5520, 5560, 5600, 5640, 5680, 5720, 5760, 5800, 5840, 5880, 5920, 5960, 6000, 6040, 6080, 6120, 6160, 6200, 6240, 6280, 6320, 6360, 6400, 6440, 6480, 6520, 6560, 6600, 6640, 6680, 6720, 6760, 6800, 6840, 6880, 6920, 6960, 7000, 7040, 7080, 7120, 7160, 7200, 7240, 7280, 7320, 7360, 7400, 7440, 7480, 7520, 7560, 7600, 7640, 7680, 7720, 7760, 7800, 7840, 7880, 7920, 7960, 8000, 8040, 8080, 8120, 8160, 8200, 8240, 8280, 8320, 8360, 8400, 8440, 8480, 8520, 8560, 8600, 8640, 8680, 8720, 8760, 8800, 8840, 8880, 8920, 8960, 9000, 9040, 9080, 9120, 9160, 9200, 9240, 9280, 9320, 9360, 9400, 9440, 9480, 9520, 9560, 9600, 9640, 9680, 9720, 9760, 9800, 9840, 9880, 9920, 9960, 10000, 10040, 10080, 10120, 10160, 10200, 
0, 41, 82, 123, 164, 205, 246, 287, 328, 369, 410, 451, 492, 533, 574, 615, 656, 697, 738, 779, 820, 861, 902, 943, 984, 1025, 1066, 1107, 1148, 1189, 1230, 1271, 1312, 1353, 1394, 1435, 1476, 1517, 1558, 1599, 1640, 1681, 1722, 1763, 1804, 1845, 1886, 1927, 1968, 2009, 2050, 2091, 2132, 2173, 2214, 2255, 2296, 2337, 2378, 2419, 2460, 2501, 2542, 2583, 2624, 2665, 2706, 2747, 2788, 2829, 2870, 2911, 2952, 2993, 3034, 3075, 3116, 3157, 3198, 3239, 3280, 3321, 3362, 3403, 3444, 3485, 3526, 3567, 3608, 3649, 3690, 3731, 3772, 3813, 3854, 3895, 3936, 3977, 4018, 4059, 4100, 4141, 4182, 4223, 4264, 4305, 4346, 4387, 4428, 4469, 4510, 4551, 4592, 4633, 4674, 4715, 4756, 4797, 4838, 4879, 4920, 4961, 5002, 5043, 5084, 5125, 5166, 5207, 5248, 5289, 5330, 5371, 5412, 5453, 5494, 5535, 5576, 5617, 5658, 5699, 5740, 5781, 5822, 5863, 5904, 5945, 5986, 6027, 6068, 6109, 6150, 6191, 6232, 6273, 6314, 6355, 6396, 6437, 6478, 6519, 6560, 6601, 6642, 6683, 6724, 6765, 6806, 6847, 6888, 6929, 6970, 7011, 7052, 7093, 7134, 7175, 7216, 7257, 7298, 7339, 7380, 7421, 7462, 7503, 7544, 7585, 7626, 7667, 7708, 7749, 7790, 7831, 7872, 7913, 7954, 7995, 8036, 8077, 8118, 8159, 8200, 8241, 8282, 8323, 8364, 8405, 8446, 8487, 8528, 8569, 8610, 8651, 8692, 8733, 8774, 8815, 8856, 8897, 8938, 8979, 9020, 9061, 9102, 9143, 9184, 9225, 9266, 9307, 9348, 9389, 9430, 9471, 9512, 9553, 9594, 9635, 9676, 9717, 9758, 9799, 9840, 9881, 9922, 9963, 10004, 10045, 10086, 10127, 10168, 10209, 10250, 10291, 10332, 10373, 10414, 10455, 
0, 42, 84, 126, 168, 210, 252, 294, 336, 378, 420, 462, 504, 546, 588, 630, 672, 714, 756, 798, 840, 882, 924, 966, 1008, 1050, 1092, 1134, 1176, 1218, 1260, 1302, 1344, 1386, 1428, 1470, 1512, 1554, 1596, 1638, 1680, 1722, 1764, 1806, 1848, 1890, 1932, 1974, 2016, 2058, 2100, 2142, 2184, 2226, 2268, 2310, 2352, 2394, 2436, 2478, 2520, 2562, 2604, 2646, 2688, 2730, 2772, 2814, 2856, 2898, 2940, 2982, 3024, 3066, 3108, 3150, 3192, 3234, 3276, 3318, 3360, 3402, 3444, 3486, 3528, 3570, 3612, 3654, 3696, 3738, 3780, 3822, 3864, 3906, 3948, 3990, 4032, 4074, 4116, 4158, 4200, 4242, 4284, 4326, 4368, 4410, 4452, 4494, 4536, 4578, 4620, 4662, 4704, 4746, 4788, 4830, 4872, 4914, 4956, 4998, 5040, 5082, 5124, 5166, 5208, 5250, 5292, 5334, 5376, 5418, 5460, 5502, 5544, 5586, 5628, 5670, 5712, 5754, 5796, 5838, 5880, 5922, 5964, 6006, 6048, 6090, 6132, 6174, 6216, 6258, 6300, 6342, 6384, 6426, 6468, 6510, 6552, 6594, 6636, 6678, 6720, 6762, 6804, 6846, 6888, 6930, 6972, 7014, 7056, 7098, 7140, 7182, 7224, 7266, 7308, 7350, 7392, 7434, 7476, 7518, 7560, 7602, 7644, 7686, 7728, 7770, 7812, 7854, 7896, 7938, 7980, 8022, 8064, 8106, 8148, 8190, 8232, 8274, 8316, 8358, 8400, 8442, 8484, 8526, 8568, 8610, 8652, 8694, 8736, 8778, 8820, 8862, 8904, 8946, 8988, 9030, 9072, 9114, 9156, 9198, 9240, 9282, 9324, 9366, 9408, 9450, 9492, 9534, 9576, 9618, 9660, 9702, 9744, 9786, 9828, 9870, 9912, 9954, 9996, 10038, 10080, 10122, 10164, 10206, 10248, 10290, 10332, 10374, 10416, 10458, 10500, 10542, 10584, 10626, 10668, 10710, 
0, 43, 86, 129, 172, 215, 258, 301, 344, 387, 430, 473, 516, 559, 602, 645, 688, 731, 774, 817, 860, 903, 946, 989, 1032, 1075, 1118, 1161, 1204, 1247, 1290, 1333, 1376, 1419, 1462, 1505, 1548, 1591, 1634, 1677, 1720, 1763, 1806, 1849, 1892, 1935, 1978, 2021, 2064, 2107, 2150, 2193, 2236, 2279, 2322, 2365, 2408, 2451, 2494, 2537, 2580, 2623, 2666, 2709, 2752, 2795, 2838, 2881, 2924, 2967, 3010, 3053, 3096, 3139, 3182, 3225, 3268, 3311, 3354, 3397, 3440, 3483, 3526, 3569, 3612, 3655, 3698, 3741, 3784, 3827, 3870, 3913, 3956, 3999, 4042, 4085, 4128, 4171, 4214, 4257, 4300, 4343, 4386, 4429, 4472, 4515, 4558, 4601, 4644, 4687, 4730, 4773, 4816, 4859, 4902, 4945, 4988, 5031, 5074, 5117, 5160, 5203, 5246, 5289, 5332, 5375, 5418, 5461, 5504, 5547, 5590, 5633, 5676, 5719, 5762, 5805, 5848, 5891, 5934, 5977, 6020, 6063, 6106, 6149, 6192, 6235, 6278, 6321, 6364, 6407, 6450, 6493, 6536, 6579, 6622, 6665, 6708, 6751, 6794, 6837, 6880, 6923, 6966, 7009, 7052, 7095, 7138, 7181, 7224, 7267, 7310, 7353, 7396, 7439, 7482, 7525, 7568, 7611, 7654, 7697, 7740, 7783, 7826, 7869, 7912, 7955, 7998, 8041, 8084, 8127, 8170, 8213, 8256, 8299, 8342, 8385, 8428, 8471, 8514, 8557, 8600, 8643, 8686, 8729, 8772, 8815, 8858, 8901, 8944, 8987, 9030, 9073, 9116, 9159, 9202, 9245, 9288, 9331, 9374, 9417, 9460, 9503, 9546, 9589, 9632, 9675, 9718, 9761, 9804, 9847, 9890, 9933, 9976, 10019, 10062, 10105, 10148, 10191, 10234, 10277, 10320, 10363, 10406, 10449, 10492, 10535, 10578, 10621, 10664, 10707, 10750, 10793, 10836, 10879, 10922, 10965, 
0, 44, 88, 132, 176, 220, 264, 308, 352, 396, 440, 484, 528, 572, 616, 660, 704, 748, 792, 836, 880, 924, 968, 1012, 1056, 1100, 1144, 1188, 1232, 1276, 1320, 1364, 1408, 1452, 1496, 1540, 1584, 1628, 1672, 1716, 1760, 1804, 1848, 1892, 1936, 1980, 2024, 2068, 2112, 2156, 2200, 2244, 2288, 2332, 2376, 2420, 2464, 2508, 2552, 2596, 2640, 2684, 2728, 2772, 2816, 2860, 2904, 2948, 2992, 3036, 3080, 3124, 3168, 3212, 3256, 3300, 3344, 3388, 3432, 3476, 3520, 3564, 3608, 3652, 3696, 3740, 3784, 3828, 3872, 3916, 3960, 4004, 4048, 4092, 4136, 4180, 4224, 4268, 4312, 4356, 4400, 4444, 4488, 4532, 4576, 4620, 4664, 4708, 4752, 4796, 4840, 4884, 4928, 4972, 5016, 5060, 5104, 5148, 5192, 5236, 5280, 5324, 5368, 5412, 5456, 5500, 5544, 5588, 5632, 5676, 5720, 5764, 5808, 5852, 5896, 5940, 5984, 6028, 6072, 6116, 6160, 6204, 6248, 6292, 6336, 6380, 6424, 6468, 6512, 6556, 6600, 6644, 6688, 6732, 6776, 6820, 6864, 6908, 6952, 6996, 7040, 7084, 7128, 7172, 7216, 7260, 7304, 7348, 7392, 7436, 7480, 7524, 7568, 7612, 7656, 7700, 7744, 7788, 7832, 7876, 7920, 7964, 8008, 8052, 8096, 8140, 8184, 8228, 8272, 8316, 8360, 8404, 8448, 8492, 8536, 8580, 8624, 8668, 8712, 8756, 8800, 8844, 8888, 8932, 8976, 9020, 9064, 9108, 9152, 9196, 9240, 9284, 9328, 9372, 9416, 9460, 9504, 9548, 9592, 9636, 9680, 9724, 9768, 9812, 9856, 9900, 9944, 9988, 10032, 10076, 10120, 10164, 10208, 10252, 10296, 10340, 10384, 10428, 10472, 10516, 10560, 10604, 10648, 10692, 10736, 10780, 10824, 10868, 10912, 10956, 11000, 11044, 11088, 11132, 11176, 11220, 
0, 45, 90, 135, 180, 225, 270, 315, 360, 405, 450, 495, 540, 585, 630, 675, 720, 765, 810, 855, 900, 945, 990, 1035, 1080, 1125, 1170, 1215, 1260, 1305, 1350, 1395, 1440, 1485, 1530, 1575, 1620, 1665, 1710, 1755, 1800, 1845, 1890, 1935, 1980, 2025, 2070, 2115, 2160, 2205, 2250, 2295, 2340, 2385, 2430, 2475, 2520, 2565, 2610, 2655, 2700, 2745, 2790, 2835, 2880, 2925, 2970, 3015, 3060, 3105, 3150, 3195, 3240, 3285, 3330, 3375, 3420, 3465, 3510, 3555, 3600, 3645, 3690, 3735, 3780, 3825, 3870, 3915, 3960, 4005, 4050, 4095, 4140, 4185, 4230, 4275, 4320, 4365, 4410, 4455, 4500, 4545, 4590, 4635, 4680, 4725, 4770, 4815, 4860, 4905, 4950, 4995, 5040, 5085, 5130, 5175, 5220, 5265, 5310, 5355, 5400, 5445, 5490, 5535, 5580, 5625, 5670, 5715, 5760, 5805, 5850, 5895, 5940, 5985, 6030, 6075, 6120, 6165, 6210, 6255, 6300, 6345, 6390, 6435, 6480, 6525, 6570, 6615, 6660, 6705, 6750, 6795, 6840, 6885, 6930, 6975, 7020, 7065, 7110, 7155, 7200, 7245, 7290, 7335, 7380, 7425, 7470, 7515, 7560, 7605, 7650, 7695, 7740, 7785, 7830, 7875, 7920, 7965, 8010, 8055, 8100, 8145, 8190, 8235, 8280, 8325, 8370, 8415, 8460, 8505, 8550, 8595, 8640, 8685, 8730, 8775, 8820, 8865, 8910, 8955, 9000, 9045, 9090, 9135, 9180, 9225, 9270, 9315, 9360, 9405, 9450, 9495, 9540, 9585, 9630, 9675, 9720, 9765, 9810, 9855, 9900, 9945, 9990, 10035, 10080, 10125, 10170, 10215, 10260, 10305, 10350, 10395, 10440, 10485, 10530, 10575, 10620, 10665, 10710, 10755, 10800, 10845, 10890, 10935, 10980, 11025, 11070, 11115, 11160, 11205, 11250, 11295, 11340, 11385, 11430, 11475, 
0, 46, 92, 138, 184, 230, 276, 322, 368, 414, 460, 506, 552, 598, 644, 690, 736, 782, 828, 874, 920, 966, 1012, 1058, 1104, 1150, 1196, 1242, 1288, 1334, 1380, 1426, 1472, 1518, 1564, 1610, 1656, 1702, 1748, 1794, 1840, 1886, 1932, 1978, 2024, 2070, 2116, 2162, 2208, 2254, 2300, 2346, 2392, 2438, 2484, 2530, 2576, 2622, 2668, 2714, 2760, 2806, 2852, 2898, 2944, 2990, 3036, 3082, 3128, 3174, 3220, 3266, 3312, 3358, 3404, 3450, 3496, 3542, 3588, 3634, 3680, 3726, 3772, 3818, 3864, 3910, 3956, 4002, 4048, 4094, 4140, 4186, 4232, 4278, 4324, 4370, 4416, 4462, 4508, 4554, 4600, 4646, 4692, 4738, 4784, 4830, 4876, 4922, 4968, 5014, 5060, 5106, 5152, 5198, 5244, 5290, 5336, 5382, 5428, 5474, 5520, 5566, 5612, 5658, 5704, 5750, 5796, 5842, 5888, 5934, 5980, 6026, 6072, 6118, 6164, 6210, 6256, 6302, 6348, 6394, 6440, 6486, 6532, 6578, 6624, 6670, 6716, 6762, 6808, 6854, 6900, 6946, 6992, 7038, 7084, 7130, 7176, 7222, 7268, 7314, 7360, 7406, 7452, 7498, 7544, 7590, 7636, 7682, 7728, 7774, 7820, 7866, 7912, 7958, 8004, 8050, 8096, 8142, 8188, 8234, 8280, 8326, 8372, 8418, 8464, 8510, 8556, 8602, 8648, 8694, 8740, 8786, 8832, 8878, 8924, 8970, 9016, 9062, 9108, 9154, 9200, 9246, 9292, 9338, 9384, 9430, 9476, 9522, 9568, 9614, 9660, 9706, 9752, 9798, 9844, 9890, 9936, 9982, 10028, 10074, 10120, 10166, 10212, 10258, 10304, 10350, 10396, 10442, 10488, 10534, 10580, 10626, 10672, 10718, 10764, 10810, 10856, 10902, 10948, 10994, 11040, 11086, 11132, 11178, 11224, 11270, 11316, 11362, 11408, 11454, 11500, 11546, 11592, 11638, 11684, 11730, 
0, 47, 94, 141, 188, 235, 282, 329, 376, 423, 470, 517, 564, 611, 658, 705, 752, 799, 846, 893, 940, 987, 1034, 1081, 1128, 1175, 1222, 1269, 1316, 1363, 1410, 1457, 1504, 1551, 1598, 1645, 1692, 1739, 1786, 1833, 1880, 1927, 1974, 2021, 2068, 2115, 2162, 2209, 2256, 2303, 2350, 2397, 2444, 2491, 2538, 2585, 2632, 2679, 2726, 2773, 2820, 2867, 2914, 2961, 3008, 3055, 3102, 3149, 3196, 3243, 3290, 3337, 3384, 3431, 3478, 3525, 3572, 3619, 3666, 3713, 3760, 3807, 3854, 3901, 3948, 3995, 4042, 4089, 4136, 4183, 4230, 4277, 4324, 4371, 4418, 4465, 4512, 4559, 4606, 4653, 4700, 4747, 4794, 4841, 4888, 4935, 4982, 5029, 5076, 5123, 5170, 5217, 5264, 5311, 5358, 5405, 5452, 5499, 5546, 5593, 5640, 5687, 5734, 5781, 5828, 5875, 5922, 5969, 6016, 6063, 6110, 6157, 6204, 6251, 6298, 6345, 6392, 6439, 6486, 6533, 6580, 6627, 6674, 6721, 6768, 6815, 6862, 6909, 6956, 7003, 7050, 7097, 7144, 7191, 7238, 7285, 7332, 7379, 7426, 7473, 7520, 7567, 7614, 7661, 7708, 7755, 7802, 7849, 7896, 7943, 7990, 8037, 8084, 8131, 8178, 8225, 8272, 8319, 8366, 8413, 8460, 8507, 8554, 8601, 8648, 8695, 8742, 8789, 8836, 8883, 8930, 8977, 9024, 9071, 9118, 9165, 9212, 9259, 9306, 9353, 9400, 9447, 9494, 9541, 9588, 9635, 9682, 9729, 9776, 9823, 9870, 9917, 9964, 10011, 10058, 10105, 10152, 10199, 10246, 10293, 10340, 10387, 10434, 10481, 10528, 10575, 10622, 10669, 10716, 10763, 10810, 10857, 10904, 10951, 10998, 11045, 11092, 11139, 11186, 11233, 11280, 11327, 11374, 11421, 11468, 11515, 11562, 11609, 11656, 11703, 11750, 11797, 11844, 11891, 11938, 11985, 
0, 48, 96, 144, 192, 240, 288, 336, 384, 432, 480, 528, 576, 624, 672, 720, 768, 816, 864, 912, 960, 1008, 1056, 1104, 1152, 1200, 1248, 1296, 1344, 1392, 1440, 1488, 1536, 1584, 1632, 1680, 1728, 1776, 1824, 1872, 1920, 1968, 2016, 2064, 2112, 2160, 2208, 2256, 2304, 2352, 2400, 2448, 2496, 2544, 2592, 2640, 2688, 2736, 2784, 2832, 2880, 2928, 2976, 3024, 3072, 3120, 3168, 3216, 3264, 3312, 3360, 3408, 3456, 3504, 3552, 3600, 3648, 3696, 3744, 3792, 3840, 3888, 3936, 3984, 4032, 4080, 4128, 4176, 4224, 4272, 4320, 4368, 4416, 4464, 4512, 4560, 4608, 4656, 4704, 4752, 4800, 4848, 4896, 4944, 4992, 5040, 5088, 5136, 5184, 5232, 5280, 5328, 5376, 5424, 5472, 5520, 5568, 5616, 5664, 5712, 5760, 5808, 5856, 5904, 5952, 6000, 6048, 6096, 6144, 6192, 6240, 6288, 6336, 6384, 6432, 6480, 6528, 6576, 6624, 6672, 6720, 6768, 6816, 6864, 6912, 6960, 7008, 7056, 7104, 7152, 7200, 7248, 7296, 7344, 7392, 7440, 7488, 7536, 7584, 7632, 7680, 7728, 7776, 7824, 7872, 7920, 7968, 8016, 8064, 8112, 8160, 8208, 8256, 8304, 8352, 8400, 8448, 8496, 8544, 8592, 8640, 8688, 8736, 8784, 8832, 8880, 8928, 8976, 9024, 9072, 9120, 9168, 9216, 9264, 9312, 9360, 9408, 9456, 9504, 9552, 9600, 9648, 9696, 9744, 9792, 9840, 9888, 9936, 9984, 10032, 10080, 10128, 10176, 10224, 10272, 10320, 10368, 10416, 10464, 10512, 10560, 10608, 10656, 10704, 10752, 10800, 10848, 10896, 10944, 10992, 11040, 11088, 11136, 11184, 11232, 11280, 11328, 11376, 11424, 11472, 11520, 11568, 11616, 11664, 11712, 11760, 11808, 11856, 11904, 11952, 12000, 12048, 12096, 12144, 12192, 12240, 
0, 49, 98, 147, 196, 245, 294, 343, 392, 441, 490, 539, 588, 637, 686, 735, 784, 833, 882, 931, 980, 1029, 1078, 1127, 1176, 1225, 1274, 1323, 1372, 1421, 1470, 1519, 1568, 1617, 1666, 1715, 1764, 1813, 1862, 1911, 1960, 2009, 2058, 2107, 2156, 2205, 2254, 2303, 2352, 2401, 2450, 2499, 2548, 2597, 2646, 2695, 2744, 2793, 2842, 2891, 2940, 2989, 3038, 3087, 3136, 3185, 3234, 3283, 3332, 3381, 3430, 3479, 3528, 3577, 3626, 3675, 3724, 3773, 3822, 3871, 3920, 3969, 4018, 4067, 4116, 4165, 4214, 4263, 4312, 4361, 4410, 4459, 4508, 4557, 4606, 4655, 4704, 4753, 4802, 4851, 4900, 4949, 4998, 5047, 5096, 5145, 5194, 5243, 5292, 5341, 5390, 5439, 5488, 5537, 5586, 5635, 5684, 5733, 5782, 5831, 5880, 5929, 5978, 6027, 6076, 6125, 6174, 6223, 6272, 6321, 6370, 6419, 6468, 6517, 6566, 6615, 6664, 6713, 6762, 6811, 6860, 6909, 6958, 7007, 7056, 7105, 7154, 7203, 7252, 7301, 7350, 7399, 7448, 7497, 7546, 7595, 7644, 7693, 7742, 7791, 7840, 7889, 7938, 7987, 8036, 8085, 8134, 8183, 8232, 8281, 8330, 8379, 8428, 8477, 8526, 8575, 8624, 8673, 8722, 8771, 8820, 8869, 8918, 8967, 9016, 9065, 9114, 9163, 9212, 9261, 9310, 9359, 9408, 9457, 9506, 9555, 9604, 9653, 9702, 9751, 9800, 9849, 9898, 9947, 9996, 10045, 10094, 10143, 10192, 10241, 10290, 10339, 10388, 10437, 10486, 10535, 10584, 10633, 10682, 10731, 10780, 10829, 10878, 10927, 10976, 11025, 11074, 11123, 11172, 11221, 11270, 11319, 11368, 11417, 11466, 11515, 11564, 11613, 11662, 11711, 11760, 11809, 11858, 11907, 11956, 12005, 12054, 12103, 12152, 12201, 12250, 12299, 12348, 12397, 12446, 12495, 
0, 50, 100, 150, 200, 250, 300, 350, 400, 450, 500, 550, 600, 650, 700, 750, 800, 850, 900, 950, 1000, 1050, 1100, 1150, 1200, 1250, 1300, 1350, 1400, 1450, 1500, 1550, 1600, 1650, 1700, 1750, 1800, 1850, 1900, 1950, 2000, 2050, 2100, 2150, 2200, 2250, 2300, 2350, 2400, 2450, 2500, 2550, 2600, 2650, 2700, 2750, 2800, 2850, 2900, 2950, 3000, 3050, 3100, 3150, 3200, 3250, 3300, 3350, 3400, 3450, 3500, 3550, 3600, 3650, 3700, 3750, 3800, 3850, 3900, 3950, 4000, 4050, 4100, 4150, 4200, 4250, 4300, 4350, 4400, 4450, 4500, 4550, 4600, 4650, 4700, 4750, 4800, 4850, 4900, 4950, 5000, 5050, 5100, 5150, 5200, 5250, 5300, 5350, 5400, 5450, 5500, 5550, 5600, 5650, 5700, 5750, 5800, 5850, 5900, 5950, 6000, 6050, 6100, 6150, 6200, 6250, 6300, 6350, 6400, 6450, 6500, 6550, 6600, 6650, 6700, 6750, 6800, 6850, 6900, 6950, 7000, 7050, 7100, 7150, 7200, 7250, 7300, 7350, 7400, 7450, 7500, 7550, 7600, 7650, 7700, 7750, 7800, 7850, 7900, 7950, 8000, 8050, 8100, 8150, 8200, 8250, 8300, 8350, 8400, 8450, 8500, 8550, 8600, 8650, 8700, 8750, 8800, 8850, 8900, 8950, 9000, 9050, 9100, 9150, 9200, 9250, 9300, 9350, 9400, 9450, 9500, 9550, 9600, 9650, 9700, 9750, 9800, 9850, 9900, 9950, 10000, 10050, 10100, 10150, 10200, 10250, 10300, 10350, 10400, 10450, 10500, 10550, 10600, 10650, 10700, 10750, 10800, 10850, 10900, 10950, 11000, 11050, 11100, 11150, 11200, 11250, 11300, 11350, 11400, 11450, 11500, 11550, 11600, 11650, 11700, 11750, 11800, 11850, 11900, 11950, 12000, 12050, 12100, 12150, 12200, 12250, 12300, 12350, 12400, 12450, 12500, 12550, 12600, 12650, 12700, 12750, 
0, 51, 102, 153, 204, 255, 306, 357, 408, 459, 510, 561, 612, 663, 714, 765, 816, 867, 918, 969, 1020, 1071, 1122, 1173, 1224, 1275, 1326, 1377, 1428, 1479, 1530, 1581, 1632, 1683, 1734, 1785, 1836, 1887, 1938, 1989, 2040, 2091, 2142, 2193, 2244, 2295, 2346, 2397, 2448, 2499, 2550, 2601, 2652, 2703, 2754, 2805, 2856, 2907, 2958, 3009, 3060, 3111, 3162, 3213, 3264, 3315, 3366, 3417, 3468, 3519, 3570, 3621, 3672, 3723, 3774, 3825, 3876, 3927, 3978, 4029, 4080, 4131, 4182, 4233, 4284, 4335, 4386, 4437, 4488, 4539, 4590, 4641, 4692, 4743, 4794, 4845, 4896, 4947, 4998, 5049, 5100, 5151, 5202, 5253, 5304, 5355, 5406, 5457, 5508, 5559, 5610, 5661, 5712, 5763, 5814, 5865, 5916, 5967, 6018, 6069, 6120, 6171, 6222, 6273, 6324, 6375, 6426, 6477, 6528, 6579, 6630, 6681, 6732, 6783, 6834, 6885, 6936, 6987, 7038, 7089, 7140, 7191, 7242, 7293, 7344, 7395, 7446, 7497, 7548, 7599, 7650, 7701, 7752, 7803, 7854, 7905, 7956, 8007, 8058, 8109, 8160, 8211, 8262, 8313, 8364, 8415, 8466, 8517, 8568, 8619, 8670, 8721, 8772, 8823, 8874, 8925, 8976, 9027, 9078, 9129, 9180, 9231, 9282, 9333, 9384, 9435, 9486, 9537, 9588, 9639, 9690, 9741, 9792, 9843, 9894, 9945, 9996, 10047, 10098, 10149, 10200, 10251, 10302, 10353, 10404, 10455, 10506, 10557, 10608, 10659, 10710, 10761, 10812, 10863, 10914, 10965, 11016, 11067, 11118, 11169, 11220, 11271, 11322, 11373, 11424, 11475, 11526, 11577, 11628, 11679, 11730, 11781, 11832, 11883, 11934, 11985, 12036, 12087, 12138, 12189, 12240, 12291, 12342, 12393, 12444, 12495, 12546, 12597, 12648, 12699, 12750, 12801, 12852, 12903, 12954, 13005, 
0, 52, 104, 156, 208, 260, 312, 364, 416, 468, 520, 572, 624, 676, 728, 780, 832, 884, 936, 988, 1040, 1092, 1144, 1196, 1248, 1300, 1352, 1404, 1456, 1508, 1560, 1612, 1664, 1716, 1768, 1820, 1872, 1924, 1976, 2028, 2080, 2132, 2184, 2236, 2288, 2340, 2392, 2444, 2496, 2548, 2600, 2652, 2704, 2756, 2808, 2860, 2912, 2964, 3016, 3068, 3120, 3172, 3224, 3276, 3328, 3380, 3432, 3484, 3536, 3588, 3640, 3692, 3744, 3796, 3848, 3900, 3952, 4004, 4056, 4108, 4160, 4212, 4264, 4316, 4368, 4420, 4472, 4524, 4576, 4628, 4680, 4732, 4784, 4836, 4888, 4940, 4992, 5044, 5096, 5148, 5200, 5252, 5304, 5356, 5408, 5460, 5512, 5564, 5616, 5668, 5720, 5772, 5824, 5876, 5928, 5980, 6032, 6084, 6136, 6188, 6240, 6292, 6344, 6396, 6448, 6500, 6552, 6604, 6656, 6708, 6760, 6812, 6864, 6916, 6968, 7020, 7072, 7124, 7176, 7228, 7280, 7332, 7384, 7436, 7488, 7540, 7592, 7644, 7696, 7748, 7800, 7852, 7904, 7956, 8008, 8060, 8112, 8164, 8216, 8268, 8320, 8372, 8424, 8476, 8528, 8580, 8632, 8684, 8736, 8788, 8840, 8892, 8944, 8996, 9048, 9100, 9152, 9204, 9256, 9308, 9360, 9412, 9464, 9516, 9568, 9620, 9672, 9724, 9776, 9828, 9880, 9932, 9984, 10036, 10088, 10140, 10192, 10244, 10296, 10348, 10400, 10452, 10504, 10556, 10608, 10660, 10712, 10764, 10816, 10868, 10920, 10972, 11024, 11076, 11128, 11180, 11232, 11284, 11336, 11388, 11440, 11492, 11544, 11596, 11648, 11700, 11752, 11804, 11856, 11908, 11960, 12012, 12064, 12116, 12168, 12220, 12272, 12324, 12376, 12428, 12480, 12532, 12584, 12636, 12688, 12740, 12792, 12844, 12896, 12948, 13000, 13052, 13104, 13156, 13208, 13260, 
0, 53, 106, 159, 212, 265, 318, 371, 424, 477, 530, 583, 636, 689, 742, 795, 848, 901, 954, 1007, 1060, 1113, 1166, 1219, 1272, 1325, 1378, 1431, 1484, 1537, 1590, 1643, 1696, 1749, 1802, 1855, 1908, 1961, 2014, 2067, 2120, 2173, 2226, 2279, 2332, 2385, 2438, 2491, 2544, 2597, 2650, 2703, 2756, 2809, 2862, 2915, 2968, 3021, 3074, 3127, 3180, 3233, 3286, 3339, 3392, 3445, 3498, 3551, 3604, 3657, 3710, 3763, 3816, 3869, 3922, 3975, 4028, 4081, 4134, 4187, 4240, 4293, 4346, 4399, 4452, 4505, 4558, 4611, 4664, 4717, 4770, 4823, 4876, 4929, 4982, 5035, 5088, 5141, 5194, 5247, 5300, 5353, 5406, 5459, 5512, 5565, 5618, 5671, 5724, 5777, 5830, 5883, 5936, 5989, 6042, 6095, 6148, 6201, 6254, 6307, 6360, 6413, 6466, 6519, 6572, 6625, 6678, 6731, 6784, 6837, 6890, 6943, 6996, 7049, 7102, 7155, 7208, 7261, 7314, 7367, 7420, 7473, 7526, 7579, 7632, 7685, 7738, 7791, 7844, 7897, 7950, 8003, 8056, 8109, 8162, 8215, 8268, 8321, 8374, 8427, 8480, 8533, 8586, 8639, 8692, 8745, 8798, 8851, 8904, 8957, 9010, 9063, 9116, 9169, 9222, 9275, 9328, 9381, 9434, 9487, 9540, 9593, 9646, 9699, 9752, 9805, 9858, 9911, 9964, 10017, 10070, 10123, 10176, 10229, 10282, 10335, 10388, 10441, 10494, 10547, 10600, 10653, 10706, 10759, 10812, 10865, 10918, 10971, 11024, 11077, 11130, 11183, 11236, 11289, 11342, 11395, 11448, 11501, 11554, 11607, 11660, 11713, 11766, 11819, 11872, 11925, 11978, 12031, 12084, 12137, 12190, 12243, 12296, 12349, 12402, 12455, 12508, 12561, 12614, 12667, 12720, 12773, 12826, 12879, 12932, 12985, 13038, 13091, 13144, 13197, 13250, 13303, 13356, 13409, 13462, 13515, 
0, 54, 108, 162, 216, 270, 324, 378, 432, 486, 540, 594, 648, 702, 756, 810, 864, 918, 972, 1026, 1080, 1134, 1188, 1242, 1296, 1350, 1404, 1458, 1512, 1566, 1620, 1674, 1728, 1782, 1836, 1890, 1944, 1998, 2052, 2106, 2160, 2214, 2268, 2322, 2376, 2430, 2484, 2538, 2592, 2646, 2700, 2754, 2808, 2862, 2916, 2970, 3024, 3078, 3132, 3186, 3240, 3294, 3348, 3402, 3456, 3510, 3564, 3618, 3672, 3726, 3780, 3834, 3888, 3942, 3996, 4050, 4104, 4158, 4212, 4266, 4320, 4374, 4428, 4482, 4536, 4590, 4644, 4698, 4752, 4806, 4860, 4914, 4968, 5022, 5076, 5130, 5184, 5238, 5292, 5346, 5400, 5454, 5508, 5562, 5616, 5670, 5724, 5778, 5832, 5886, 5940, 5994, 6048, 6102, 6156, 6210, 6264, 6318, 6372, 6426, 6480, 6534, 6588, 6642, 6696, 6750, 6804, 6858, 6912, 6966, 7020, 7074, 7128, 7182, 7236, 7290, 7344, 7398, 7452, 7506, 7560, 7614, 7668, 7722, 7776, 7830, 7884, 7938, 7992, 8046, 8100, 8154, 8208, 8262, 8316, 8370, 8424, 8478, 8532, 8586, 8640, 8694, 8748, 8802, 8856, 8910, 8964, 9018, 9072, 9126, 9180, 9234, 9288, 9342, 9396, 9450, 9504, 9558, 9612, 9666, 9720, 9774, 9828, 9882, 9936, 9990, 10044, 10098, 10152, 10206, 10260, 10314, 10368, 10422, 10476, 10530, 10584, 10638, 10692, 10746, 10800, 10854, 10908, 10962, 11016, 11070, 11124, 11178, 11232, 11286, 11340, 11394, 11448, 11502, 11556, 11610, 11664, 11718, 11772, 11826, 11880, 11934, 11988, 12042, 12096, 12150, 12204, 12258, 12312, 12366, 12420, 12474, 12528, 12582, 12636, 12690, 12744, 12798, 12852, 12906, 12960, 13014, 13068, 13122, 13176, 13230, 13284, 13338, 13392, 13446, 13500, 13554, 13608, 13662, 13716, 13770, 
0, 55, 110, 165, 220, 275, 330, 385, 440, 495, 550, 605, 660, 715, 770, 825, 880, 935, 990, 1045, 1100, 1155, 1210, 1265, 1320, 1375, 1430, 1485, 1540, 1595, 1650, 1705, 1760, 1815, 1870, 1925, 1980, 2035, 2090, 2145, 2200, 2255, 2310, 2365, 2420, 2475, 2530, 2585, 2640, 2695, 2750, 2805, 2860, 2915, 2970, 3025, 3080, 3135, 3190, 3245, 3300, 3355, 3410, 3465, 3520, 3575, 3630, 3685, 3740, 3795, 3850, 3905, 3960, 4015, 4070, 4125, 4180, 4235, 4290, 4345, 4400, 4455, 4510, 4565, 4620, 4675, 4730, 4785, 4840, 4895, 4950, 5005, 5060, 5115, 5170, 5225, 5280, 5335, 5390, 5445, 5500, 5555, 5610, 5665, 5720, 5775, 5830, 5885, 5940, 5995, 6050, 6105, 6160, 6215, 6270, 6325, 6380, 6435, 6490, 6545, 6600, 6655, 6710, 6765, 6820, 6875, 6930, 6985, 7040, 7095, 7150, 7205, 7260, 7315, 7370, 7425, 7480, 7535, 7590, 7645, 7700, 7755, 7810, 7865, 7920, 7975, 8030, 8085, 8140, 8195, 8250, 8305, 8360, 8415, 8470, 8525, 8580, 8635, 8690, 8745, 8800, 8855, 8910, 8965, 9020, 9075, 9130, 9185, 9240, 9295, 9350, 9405, 9460, 9515, 9570, 9625, 9680, 9735, 9790, 9845, 9900, 9955, 10010, 10065, 10120, 10175, 10230, 10285, 10340, 10395, 10450, 10505, 10560, 10615, 10670, 10725, 10780, 10835, 10890, 10945, 11000, 11055, 11110, 11165, 11220, 11275, 11330, 11385, 11440, 11495, 11550, 11605, 11660, 11715, 11770, 11825, 11880, 11935, 11990, 12045, 12100, 12155, 12210, 12265, 12320, 12375, 12430, 12485, 12540, 12595, 12650, 12705, 12760, 12815, 12870, 12925, 12980, 13035, 13090, 13145, 13200, 13255, 13310, 13365, 13420, 13475, 13530, 13585, 13640, 13695, 13750, 13805, 13860, 13915, 13970, 14025, 
0, 56, 112, 168, 224, 280, 336, 392, 448, 504, 560, 616, 672, 728, 784, 840, 896, 952, 1008, 1064, 1120, 1176, 1232, 1288, 1344, 1400, 1456, 1512, 1568, 1624, 1680, 1736, 1792, 1848, 1904, 1960, 2016, 2072, 2128, 2184, 2240, 2296, 2352, 2408, 2464, 2520, 2576, 2632, 2688, 2744, 2800, 2856, 2912, 2968, 3024, 3080, 3136, 3192, 3248, 3304, 3360, 3416, 3472, 3528, 3584, 3640, 3696, 3752, 3808, 3864, 3920, 3976, 4032, 4088, 4144, 4200, 4256, 4312, 4368, 4424, 4480, 4536, 4592, 4648, 4704, 4760, 4816, 4872, 4928, 4984, 5040, 5096, 5152, 5208, 5264, 5320, 5376, 5432, 5488, 5544, 5600, 5656, 5712, 5768, 5824, 5880, 5936, 5992, 6048, 6104, 6160, 6216, 6272, 6328, 6384, 6440, 6496, 6552, 6608, 6664, 6720, 6776, 6832, 6888, 6944, 7000, 7056, 7112, 7168, 7224, 7280, 7336, 7392, 7448, 7504, 7560, 7616, 7672, 7728, 7784, 7840, 7896, 7952, 8008, 8064, 8120, 8176, 8232, 8288, 8344, 8400, 8456, 8512, 8568, 8624, 8680, 8736, 8792, 8848, 8904, 8960, 9016, 9072, 9128, 9184, 9240, 9296, 9352, 9408, 9464, 9520, 9576, 9632, 9688, 9744, 9800, 9856, 9912, 9968, 10024, 10080, 10136, 10192, 10248, 10304, 10360, 10416, 10472, 10528, 10584, 10640, 10696, 10752, 10808, 10864, 10920, 10976, 11032, 11088, 11144, 11200, 11256, 11312, 11368, 11424, 11480, 11536, 11592, 11648, 11704, 11760, 11816, 11872, 11928, 11984, 12040, 12096, 12152, 12208, 12264, 12320, 12376, 12432, 12488, 12544, 12600, 12656, 12712, 12768, 12824, 12880, 12936, 12992, 13048, 13104, 13160, 13216, 13272, 13328, 13384, 13440, 13496, 13552, 13608, 13664, 13720, 13776, 13832, 13888, 13944, 14000, 14056, 14112, 14168, 14224, 14280, 
0, 57, 114, 171, 228, 285, 342, 399, 456, 513, 570, 627, 684, 741, 798, 855, 912, 969, 1026, 1083, 1140, 1197, 1254, 1311, 1368, 1425, 1482, 1539, 1596, 1653, 1710, 1767, 1824, 1881, 1938, 1995, 2052, 2109, 2166, 2223, 2280, 2337, 2394, 2451, 2508, 2565, 2622, 2679, 2736, 2793, 2850, 2907, 2964, 3021, 3078, 3135, 3192, 3249, 3306, 3363, 3420, 3477, 3534, 3591, 3648, 3705, 3762, 3819, 3876, 3933, 3990, 4047, 4104, 4161, 4218, 4275, 4332, 4389, 4446, 4503, 4560, 4617, 4674, 4731, 4788, 4845, 4902, 4959, 5016, 5073, 5130, 5187, 5244, 5301, 5358, 5415, 5472, 5529, 5586, 5643, 5700, 5757, 5814, 5871, 5928, 5985, 6042, 6099, 6156, 6213, 6270, 6327, 6384, 6441, 6498, 6555, 6612, 6669, 6726, 6783, 6840, 6897, 6954, 7011, 7068, 7125, 7182, 7239, 7296, 7353, 7410, 7467, 7524, 7581, 7638, 7695, 7752, 7809, 7866, 7923, 7980, 8037, 8094, 8151, 8208, 8265, 8322, 8379, 8436, 8493, 8550, 8607, 8664, 8721, 8778, 8835, 8892, 8949, 9006, 9063, 9120, 9177, 9234, 9291, 9348, 9405, 9462, 9519, 9576, 9633, 9690, 9747, 9804, 9861, 9918, 9975, 10032, 10089, 10146, 10203, 10260, 10317, 10374, 10431, 10488, 10545, 10602, 10659, 10716, 10773, 10830, 10887, 10944, 11001, 11058, 11115, 11172, 11229, 11286, 11343, 11400, 11457, 11514, 11571, 11628, 11685, 11742, 11799, 11856, 11913, 11970, 12027, 12084, 12141, 12198, 12255, 12312, 12369, 12426, 12483, 12540, 12597, 12654, 12711, 12768, 12825, 12882, 12939, 12996, 13053, 13110, 13167, 13224, 13281, 13338, 13395, 13452, 13509, 13566, 13623, 13680, 13737, 13794, 13851, 13908, 13965, 14022, 14079, 14136, 14193, 14250, 14307, 14364, 14421, 14478, 14535, 
0, 58, 116, 174, 232, 290, 348, 406, 464, 522, 580, 638, 696, 754, 812, 870, 928, 986, 1044, 1102, 1160, 1218, 1276, 1334, 1392, 1450, 1508, 1566, 1624, 1682, 1740, 1798, 1856, 1914, 1972, 2030, 2088, 2146, 2204, 2262, 2320, 2378, 2436, 2494, 2552, 2610, 2668, 2726, 2784, 2842, 2900, 2958, 3016, 3074, 3132, 3190, 3248, 3306, 3364, 3422, 3480, 3538, 3596, 3654, 3712, 3770, 3828, 3886, 3944, 4002, 4060, 4118, 4176, 4234, 4292, 4350, 4408, 4466, 4524, 4582, 4640, 4698, 4756, 4814, 4872, 4930, 4988, 5046, 5104, 5162, 5220, 5278, 5336, 5394, 5452, 5510, 5568, 5626, 5684, 5742, 5800, 5858, 5916, 5974, 6032, 6090, 6148, 6206, 6264, 6322, 6380, 6438, 6496, 6554, 6612, 6670, 6728, 6786, 6844, 6902, 6960, 7018, 7076, 7134, 7192, 7250, 7308, 7366, 7424, 7482, 7540, 7598, 7656, 7714, 7772, 7830, 7888, 7946, 8004, 8062, 8120, 8178, 8236, 8294, 8352, 8410, 8468, 8526, 8584, 8642, 8700, 8758, 8816, 8874, 8932, 8990, 9048, 9106, 9164, 9222, 9280, 9338, 9396, 9454, 9512, 9570, 9628, 9686, 9744, 9802, 9860, 9918, 9976, 10034, 10092, 10150, 10208, 10266, 10324, 10382, 10440, 10498, 10556, 10614, 10672, 10730, 10788, 10846, 10904, 10962, 11020, 11078, 11136, 11194, 11252, 11310, 11368, 11426, 11484, 11542, 11600, 11658, 11716, 11774, 11832, 11890, 11948, 12006, 12064, 12122, 12180, 12238, 12296, 12354, 12412, 12470, 12528, 12586, 12644, 12702, 12760, 12818, 12876, 12934, 12992, 13050, 13108, 13166, 13224, 13282, 13340, 13398, 13456, 13514, 13572, 13630, 13688, 13746, 13804, 13862, 13920, 13978, 14036, 14094, 14152, 14210, 14268, 14326, 14384, 14442, 14500, 14558, 14616, 14674, 14732, 14790, 
0, 59, 118, 177, 236, 295, 354, 413, 472, 531, 590, 649, 708, 767, 826, 885, 944, 1003, 1062, 1121, 1180, 1239, 1298, 1357, 1416, 1475, 1534, 1593, 1652, 1711, 1770, 1829, 1888, 1947, 2006, 2065, 2124, 2183, 2242, 2301, 2360, 2419, 2478, 2537, 2596, 2655, 2714, 2773, 2832, 2891, 2950, 3009, 3068, 3127, 3186, 3245, 3304, 3363, 3422, 3481, 3540, 3599, 3658, 3717, 3776, 3835, 3894, 3953, 4012, 4071, 4130, 4189, 4248, 4307, 4366, 4425, 4484, 4543, 4602, 4661, 4720, 4779, 4838, 4897, 4956, 5015, 5074, 5133, 5192, 5251, 5310, 5369, 5428, 5487, 5546, 5605, 5664, 5723, 5782, 5841, 5900, 5959, 6018, 6077, 6136, 6195, 6254, 6313, 6372, 6431, 6490, 6549, 6608, 6667, 6726, 6785, 6844, 6903, 6962, 7021, 7080, 7139, 7198, 7257, 7316, 7375, 7434, 7493, 7552, 7611, 7670, 7729, 7788, 7847, 7906, 7965, 8024, 8083, 8142, 8201, 8260, 8319, 8378, 8437, 8496, 8555, 8614, 8673, 8732, 8791, 8850, 8909, 8968, 9027, 9086, 9145, 9204, 9263, 9322, 9381, 9440, 9499, 9558, 9617, 9676, 9735, 9794, 9853, 9912, 9971, 10030, 10089, 10148, 10207, 10266, 10325, 10384, 10443, 10502, 10561, 10620, 10679, 10738, 10797, 10856, 10915, 10974, 11033, 11092, 11151, 11210, 11269, 11328, 11387, 11446, 11505, 11564, 11623, 11682, 11741, 11800, 11859, 11918, 11977, 12036, 12095, 12154, 12213, 12272, 12331, 12390, 12449, 12508, 12567, 12626, 12685, 12744, 12803, 12862, 12921, 12980, 13039, 13098, 13157, 13216, 13275, 13334, 13393, 13452, 13511, 13570, 13629, 13688, 13747, 13806, 13865, 13924, 13983, 14042, 14101, 14160, 14219, 14278, 14337, 14396, 14455, 14514, 14573, 14632, 14691, 14750, 14809, 14868, 14927, 14986, 15045, 
0, 60, 120, 180, 240, 300, 360, 420, 480, 540, 600, 660, 720, 780, 840, 900, 960, 1020, 1080, 1140, 1200, 1260, 1320, 1380, 1440, 1500, 1560, 1620, 1680, 1740, 1800, 1860, 1920, 1980, 2040, 2100, 2160, 2220, 2280, 2340, 2400, 2460, 2520, 2580, 2640, 2700, 2760, 2820, 2880, 2940, 3000, 3060, 3120, 3180, 3240, 3300, 3360, 3420, 3480, 3540, 3600, 3660, 3720, 3780, 3840, 3900, 3960, 4020, 4080, 4140, 4200, 4260, 4320, 4380, 4440, 4500, 4560, 4620, 4680, 4740, 4800, 4860, 4920, 4980, 5040, 5100, 5160, 5220, 5280, 5340, 5400, 5460, 5520, 5580, 5640, 5700, 5760, 5820, 5880, 5940, 6000, 6060, 6120, 6180, 6240, 6300, 6360, 6420, 6480, 6540, 6600, 6660, 6720, 6780, 6840, 6900, 6960, 7020, 7080, 7140, 7200, 7260, 7320, 7380, 7440, 7500, 7560, 7620, 7680, 7740, 7800, 7860, 7920, 7980, 8040, 8100, 8160, 8220, 8280, 8340, 8400, 8460, 8520, 8580, 8640, 8700, 8760, 8820, 8880, 8940, 9000, 9060, 9120, 9180, 9240, 9300, 9360, 9420, 9480, 9540, 9600, 9660, 9720, 9780, 9840, 9900, 9960, 10020, 10080, 10140, 10200, 10260, 10320, 10380, 10440, 10500, 10560, 10620, 10680, 10740, 10800, 10860, 10920, 10980, 11040, 11100, 11160, 11220, 11280, 11340, 11400, 11460, 11520, 11580, 11640, 11700, 11760, 11820, 11880, 11940, 12000, 12060, 12120, 12180, 12240, 12300, 12360, 12420, 12480, 12540, 12600, 12660, 12720, 12780, 12840, 12900, 12960, 13020, 13080, 13140, 13200, 13260, 13320, 13380, 13440, 13500, 13560, 13620, 13680, 13740, 13800, 13860, 13920, 13980, 14040, 14100, 14160, 14220, 14280, 14340, 14400, 14460, 14520, 14580, 14640, 14700, 14760, 14820, 14880, 14940, 15000, 15060, 15120, 15180, 15240, 15300, 
0, 61, 122, 183, 244, 305, 366, 427, 488, 549, 610, 671, 732, 793, 854, 915, 976, 1037, 1098, 1159, 1220, 1281, 1342, 1403, 1464, 1525, 1586, 1647, 1708, 1769, 1830, 1891, 1952, 2013, 2074, 2135, 2196, 2257, 2318, 2379, 2440, 2501, 2562, 2623, 2684, 2745, 2806, 2867, 2928, 2989, 3050, 3111, 3172, 3233, 3294, 3355, 3416, 3477, 3538, 3599, 3660, 3721, 3782, 3843, 3904, 3965, 4026, 4087, 4148, 4209, 4270, 4331, 4392, 4453, 4514, 4575, 4636, 4697, 4758, 4819, 4880, 4941, 5002, 5063, 5124, 5185, 5246, 5307, 5368, 5429, 5490, 5551, 5612, 5673, 5734, 5795, 5856, 5917, 5978, 6039, 6100, 6161, 6222, 6283, 6344, 6405, 6466, 6527, 6588, 6649, 6710, 6771, 6832, 6893, 6954, 7015, 7076, 7137, 7198, 7259, 7320, 7381, 7442, 7503, 7564, 7625, 7686, 7747, 7808, 7869, 7930, 7991, 8052, 8113, 8174, 8235, 8296, 8357, 8418, 8479, 8540, 8601, 8662, 8723, 8784, 8845, 8906, 8967, 9028, 9089, 9150, 9211, 9272, 9333, 9394, 9455, 9516, 9577, 9638, 9699, 9760, 9821, 9882, 9943, 10004, 10065, 10126, 10187, 10248, 10309, 10370, 10431, 10492, 10553, 10614, 10675, 10736, 10797, 10858, 10919, 10980, 11041, 11102, 11163, 11224, 11285, 11346, 11407, 11468, 11529, 11590, 11651, 11712, 11773, 11834, 11895, 11956, 12017, 12078, 12139, 12200, 12261, 12322, 12383, 12444, 12505, 12566, 12627, 12688, 12749, 12810, 12871, 12932, 12993, 13054, 13115, 13176, 13237, 13298, 13359, 13420, 13481, 13542, 13603, 13664, 13725, 13786, 13847, 13908, 13969, 14030, 14091, 14152, 14213, 14274, 14335, 14396, 14457, 14518, 14579, 14640, 14701, 14762, 14823, 14884, 14945, 15006, 15067, 15128, 15189, 15250, 15311, 15372, 15433, 15494, 15555, 
0, 62, 124, 186, 248, 310, 372, 434, 496, 558, 620, 682, 744, 806, 868, 930, 992, 1054, 1116, 1178, 1240, 1302, 1364, 1426, 1488, 1550, 1612, 1674, 1736, 1798, 1860, 1922, 1984, 2046, 2108, 2170, 2232, 2294, 2356, 2418, 2480, 2542, 2604, 2666, 2728, 2790, 2852, 2914, 2976, 3038, 3100, 3162, 3224, 3286, 3348, 3410, 3472, 3534, 3596, 3658, 3720, 3782, 3844, 3906, 3968, 4030, 4092, 4154, 4216, 4278, 4340, 4402, 4464, 4526, 4588, 4650, 4712, 4774, 4836, 4898, 4960, 5022, 5084, 5146, 5208, 5270, 5332, 5394, 5456, 5518, 5580, 5642, 5704, 5766, 5828, 5890, 5952, 6014, 6076, 6138, 6200, 6262, 6324, 6386, 6448, 6510, 6572, 6634, 6696, 6758, 6820, 6882, 6944, 7006, 7068, 7130, 7192, 7254, 7316, 7378, 7440, 7502, 7564, 7626, 7688, 7750, 7812, 7874, 7936, 7998, 8060, 8122, 8184, 8246, 8308, 8370, 8432, 8494, 8556, 8618, 8680, 8742, 8804, 8866, 8928, 8990, 9052, 9114, 9176, 9238, 9300, 9362, 9424, 9486, 9548, 9610, 9672, 9734, 9796, 9858, 9920, 9982, 10044, 10106, 10168, 10230, 10292, 10354, 10416, 10478, 10540, 10602, 10664, 10726, 10788, 10850, 10912, 10974, 11036, 11098, 11160, 11222, 11284, 11346, 11408, 11470, 11532, 11594, 11656, 11718, 11780, 11842, 11904, 11966, 12028, 12090, 12152, 12214, 12276, 12338, 12400, 12462, 12524, 12586, 12648, 12710, 12772, 12834, 12896, 12958, 13020, 13082, 13144, 13206, 13268, 13330, 13392, 13454, 13516, 13578, 13640, 13702, 13764, 13826, 13888, 13950, 14012, 14074, 14136, 14198, 14260, 14322, 14384, 14446, 14508, 14570, 14632, 14694, 14756, 14818, 14880, 14942, 15004, 15066, 15128, 15190, 15252, 15314, 15376, 15438, 15500, 15562, 15624, 15686, 15748, 15810, 
0, 63, 126, 189, 252, 315, 378, 441, 504, 567, 630, 693, 756, 819, 882, 945, 1008, 1071, 1134, 1197, 1260, 1323, 1386, 1449, 1512, 1575, 1638, 1701, 1764, 1827, 1890, 1953, 2016, 2079, 2142, 2205, 2268, 2331, 2394, 2457, 2520, 2583, 2646, 2709, 2772, 2835, 2898, 2961, 3024, 3087, 3150, 3213, 3276, 3339, 3402, 3465, 3528, 3591, 3654, 3717, 3780, 3843, 3906, 3969, 4032, 4095, 4158, 4221, 4284, 4347, 4410, 4473, 4536, 4599, 4662, 4725, 4788, 4851, 4914, 4977, 5040, 5103, 5166, 5229, 5292, 5355, 5418, 5481, 5544, 5607, 5670, 5733, 5796, 5859, 5922, 5985, 6048, 6111, 6174, 6237, 6300, 6363, 6426, 6489, 6552, 6615, 6678, 6741, 6804, 6867, 6930, 6993, 7056, 7119, 7182, 7245, 7308, 7371, 7434, 7497, 7560, 7623, 7686, 7749, 7812, 7875, 7938, 8001, 8064, 8127, 8190, 8253, 8316, 8379, 8442, 8505, 8568, 8631, 8694, 8757, 8820, 8883, 8946, 9009, 9072, 9135, 9198, 9261, 9324, 9387, 9450, 9513, 9576, 9639, 9702, 9765, 9828, 9891, 9954, 10017, 10080, 10143, 10206, 10269, 10332, 10395, 10458, 10521, 10584, 10647, 10710, 10773, 10836, 10899, 10962, 11025, 11088, 11151, 11214, 11277, 11340, 11403, 11466, 11529, 11592, 11655, 11718, 11781, 11844, 11907, 11970, 12033, 12096, 12159, 12222, 12285, 12348, 12411, 12474, 12537, 12600, 12663, 12726, 12789, 12852, 12915, 12978, 13041, 13104, 13167, 13230, 13293, 13356, 13419, 13482, 13545, 13608, 13671, 13734, 13797, 13860, 13923, 13986, 14049, 14112, 14175, 14238, 14301, 14364, 14427, 14490, 14553, 14616, 14679, 14742, 14805, 14868, 14931, 14994, 15057, 15120, 15183, 15246, 15309, 15372, 15435, 15498, 15561, 15624, 15687, 15750, 15813, 15876, 15939, 16002, 16065, 
0, 64, 128, 192, 256, 320, 384, 448, 512, 576, 640, 704, 768, 832, 896, 960, 1024, 1088, 1152, 1216, 1280, 1344, 1408, 1472, 1536, 1600, 1664, 1728, 1792, 1856, 1920, 1984, 2048, 2112, 2176, 2240, 2304, 2368, 2432, 2496, 2560, 2624, 2688, 2752, 2816, 2880, 2944, 3008, 3072, 3136, 3200, 3264, 3328, 3392, 3456, 3520, 3584, 3648, 3712, 3776, 3840, 3904, 3968, 4032, 4096, 4160, 4224, 4288, 4352, 4416, 4480, 4544, 4608, 4672, 4736, 4800, 4864, 4928, 4992, 5056, 5120, 5184, 5248, 5312, 5376, 5440, 5504, 5568, 5632, 5696, 5760, 5824, 5888, 5952, 6016, 6080, 6144, 6208, 6272, 6336, 6400, 6464, 6528, 6592, 6656, 6720, 6784, 6848, 6912, 6976, 7040, 7104, 7168, 7232, 7296, 7360, 7424, 7488, 7552, 7616, 7680, 7744, 7808, 7872, 7936, 8000, 8064, 8128, 8192, 8256, 8320, 8384, 8448, 8512, 8576, 8640, 8704, 8768, 8832, 8896, 8960, 9024, 9088, 9152, 9216, 9280, 9344, 9408, 9472, 9536, 9600, 9664, 9728, 9792, 9856, 9920, 9984, 10048, 10112, 10176, 10240, 10304, 10368, 10432, 10496, 10560, 10624, 10688, 10752, 10816, 10880, 10944, 11008, 11072, 11136, 11200, 11264, 11328, 11392, 11456, 11520, 11584, 11648, 11712, 11776, 11840, 11904, 11968, 12032, 12096, 12160, 12224, 12288, 12352, 12416, 12480, 12544, 12608, 12672, 12736, 12800, 12864, 12928, 12992, 13056, 13120, 13184, 13248, 13312, 13376, 13440, 13504, 13568, 13632, 13696, 13760, 13824, 13888, 13952, 14016, 14080, 14144, 14208, 14272, 14336, 14400, 14464, 14528, 14592, 14656, 14720, 14784, 14848, 14912, 14976, 15040, 15104, 15168, 15232, 15296, 15360, 15424, 15488, 15552, 15616, 15680, 15744, 15808, 15872, 15936, 16000, 16064, 16128, 16192, 16256, 16320, 
0, 65, 130, 195, 260, 325, 390, 455, 520, 585, 650, 715, 780, 845, 910, 975, 1040, 1105, 1170, 1235, 1300, 1365, 1430, 1495, 1560, 1625, 1690, 1755, 1820, 1885, 1950, 2015, 2080, 2145, 2210, 2275, 2340, 2405, 2470, 2535, 2600, 2665, 2730, 2795, 2860, 2925, 2990, 3055, 3120, 3185, 3250, 3315, 3380, 3445, 3510, 3575, 3640, 3705, 3770, 3835, 3900, 3965, 4030, 4095, 4160, 4225, 4290, 4355, 4420, 4485, 4550, 4615, 4680, 4745, 4810, 4875, 4940, 5005, 5070, 5135, 5200, 5265, 5330, 5395, 5460, 5525, 5590, 5655, 5720, 5785, 5850, 5915, 5980, 6045, 6110, 6175, 6240, 6305, 6370, 6435, 6500, 6565, 6630, 6695, 6760, 6825, 6890, 6955, 7020, 7085, 7150, 7215, 7280, 7345, 7410, 7475, 7540, 7605, 7670, 7735, 7800, 7865, 7930, 7995, 8060, 8125, 8190, 8255, 8320, 8385, 8450, 8515, 8580, 8645, 8710, 8775, 8840, 8905, 8970, 9035, 9100, 9165, 9230, 9295, 9360, 9425, 9490, 9555, 9620, 9685, 9750, 9815, 9880, 9945, 10010, 10075, 10140, 10205, 10270, 10335, 10400, 10465, 10530, 10595, 10660, 10725, 10790, 10855, 10920, 10985, 11050, 11115, 11180, 11245, 11310, 11375, 11440, 11505, 11570, 11635, 11700, 11765, 11830, 11895, 11960, 12025, 12090, 12155, 12220, 12285, 12350, 12415, 12480, 12545, 12610, 12675, 12740, 12805, 12870, 12935, 13000, 13065, 13130, 13195, 13260, 13325, 13390, 13455, 13520, 13585, 13650, 13715, 13780, 13845, 13910, 13975, 14040, 14105, 14170, 14235, 14300, 14365, 14430, 14495, 14560, 14625, 14690, 14755, 14820, 14885, 14950, 15015, 15080, 15145, 15210, 15275, 15340, 15405, 15470, 15535, 15600, 15665, 15730, 15795, 15860, 15925, 15990, 16055, 16120, 16185, 16250, 16315, 16380, 16445, 16510, 16575, 
0, 66, 132, 198, 264, 330, 396, 462, 528, 594, 660, 726, 792, 858, 924, 990, 1056, 1122, 1188, 1254, 1320, 1386, 1452, 1518, 1584, 1650, 1716, 1782, 1848, 1914, 1980, 2046, 2112, 2178, 2244, 2310, 2376, 2442, 2508, 2574, 2640, 2706, 2772, 2838, 2904, 2970, 3036, 3102, 3168, 3234, 3300, 3366, 3432, 3498, 3564, 3630, 3696, 3762, 3828, 3894, 3960, 4026, 4092, 4158, 4224, 4290, 4356, 4422, 4488, 4554, 4620, 4686, 4752, 4818, 4884, 4950, 5016, 5082, 5148, 5214, 5280, 5346, 5412, 5478, 5544, 5610, 5676, 5742, 5808, 5874, 5940, 6006, 6072, 6138, 6204, 6270, 6336, 6402, 6468, 6534, 6600, 6666, 6732, 6798, 6864, 6930, 6996, 7062, 7128, 7194, 7260, 7326, 7392, 7458, 7524, 7590, 7656, 7722, 7788, 7854, 7920, 7986, 8052, 8118, 8184, 8250, 8316, 8382, 8448, 8514, 8580, 8646, 8712, 8778, 8844, 8910, 8976, 9042, 9108, 9174, 9240, 9306, 9372, 9438, 9504, 9570, 9636, 9702, 9768, 9834, 9900, 9966, 10032, 10098, 10164, 10230, 10296, 10362, 10428, 10494, 10560, 10626, 10692, 10758, 10824, 10890, 10956, 11022, 11088, 11154, 11220, 11286, 11352, 11418, 11484, 11550, 11616, 11682, 11748, 11814, 11880, 11946, 12012, 12078, 12144, 12210, 12276, 12342, 12408, 12474, 12540, 12606, 12672, 12738, 12804, 12870, 12936, 13002, 13068, 13134, 13200, 13266, 13332, 13398, 13464, 13530, 13596, 13662, 13728, 13794, 13860, 13926, 13992, 14058, 14124, 14190, 14256, 14322, 14388, 14454, 14520, 14586, 14652, 14718, 14784, 14850, 14916, 14982, 15048, 15114, 15180, 15246, 15312, 15378, 15444, 15510, 15576, 15642, 15708, 15774, 15840, 15906, 15972, 16038, 16104, 16170, 16236, 16302, 16368, 16434, 16500, 16566, 16632, 16698, 16764, 16830, 
0, 67, 134, 201, 268, 335, 402, 469, 536, 603, 670, 737, 804, 871, 938, 1005, 1072, 1139, 1206, 1273, 1340, 1407, 1474, 1541, 1608, 1675, 1742, 1809, 1876, 1943, 2010, 2077, 2144, 2211, 2278, 2345, 2412, 2479, 2546, 2613, 2680, 2747, 2814, 2881, 2948, 3015, 3082, 3149, 3216, 3283, 3350, 3417, 3484, 3551, 3618, 3685, 3752, 3819, 3886, 3953, 4020, 4087, 4154, 4221, 4288, 4355, 4422, 4489, 4556, 4623, 4690, 4757, 4824, 4891, 4958, 5025, 5092, 5159, 5226, 5293, 5360, 5427, 5494, 5561, 5628, 5695, 5762, 5829, 5896, 5963, 6030, 6097, 6164, 6231, 6298, 6365, 6432, 6499, 6566, 6633, 6700, 6767, 6834, 6901, 6968, 7035, 7102, 7169, 7236, 7303, 7370, 7437, 7504, 7571, 7638, 7705, 7772, 7839, 7906, 7973, 8040, 8107, 8174, 8241, 8308, 8375, 8442, 8509, 8576, 8643, 8710, 8777, 8844, 8911, 8978, 9045, 9112, 9179, 9246, 9313, 9380, 9447, 9514, 9581, 9648, 9715, 9782, 9849, 9916, 9983, 10050, 10117, 10184, 10251, 10318, 10385, 10452, 10519, 10586, 10653, 10720, 10787, 10854, 10921, 10988, 11055, 11122, 11189, 11256, 11323, 11390, 11457, 11524, 11591, 11658, 11725, 11792, 11859, 11926, 11993, 12060, 12127, 12194, 12261, 12328, 12395, 12462, 12529, 12596, 12663, 12730, 12797, 12864, 12931, 12998, 13065, 13132, 13199, 13266, 13333, 13400, 13467, 13534, 13601, 13668, 13735, 13802, 13869, 13936, 14003, 14070, 14137, 14204, 14271, 14338, 14405, 14472, 14539, 14606, 14673, 14740, 14807, 14874, 14941, 15008, 15075, 15142, 15209, 15276, 15343, 15410, 15477, 15544, 15611, 15678, 15745, 15812, 15879, 15946, 16013, 16080, 16147, 16214, 16281, 16348, 16415, 16482, 16549, 16616, 16683, 16750, 16817, 16884, 16951, 17018, 17085, 
0, 68, 136, 204, 272, 340, 408, 476, 544, 612, 680, 748, 816, 884, 952, 1020, 1088, 1156, 1224, 1292, 1360, 1428, 1496, 1564, 1632, 1700, 1768, 1836, 1904, 1972, 2040, 2108, 2176, 2244, 2312, 2380, 2448, 2516, 2584, 2652, 2720, 2788, 2856, 2924, 2992, 3060, 3128, 3196, 3264, 3332, 3400, 3468, 3536, 3604, 3672, 3740, 3808, 3876, 3944, 4012, 4080, 4148, 4216, 4284, 4352, 4420, 4488, 4556, 4624, 4692, 4760, 4828, 4896, 4964, 5032, 5100, 5168, 5236, 5304, 5372, 5440, 5508, 5576, 5644, 5712, 5780, 5848, 5916, 5984, 6052, 6120, 6188, 6256, 6324, 6392, 6460, 6528, 6596, 6664, 6732, 6800, 6868, 6936, 7004, 7072, 7140, 7208, 7276, 7344, 7412, 7480, 7548, 7616, 7684, 7752, 7820, 7888, 7956, 8024, 8092, 8160, 8228, 8296, 8364, 8432, 8500, 8568, 8636, 8704, 8772, 8840, 8908, 8976, 9044, 9112, 9180, 9248, 9316, 9384, 9452, 9520, 9588, 9656, 9724, 9792, 9860, 9928, 9996, 10064, 10132, 10200, 10268, 10336, 10404, 10472, 10540, 10608, 10676, 10744, 10812, 10880, 10948, 11016, 11084, 11152, 11220, 11288, 11356, 11424, 11492, 11560, 11628, 11696, 11764, 11832, 11900, 11968, 12036, 12104, 12172, 12240, 12308, 12376, 12444, 12512, 12580, 12648, 12716, 12784, 12852, 12920, 12988, 13056, 13124, 13192, 13260, 13328, 13396, 13464, 13532, 13600, 13668, 13736, 13804, 13872, 13940, 14008, 14076, 14144, 14212, 14280, 14348, 14416, 14484, 14552, 14620, 14688, 14756, 14824, 14892, 14960, 15028, 15096, 15164, 15232, 15300, 15368, 15436, 15504, 15572, 15640, 15708, 15776, 15844, 15912, 15980, 16048, 16116, 16184, 16252, 16320, 16388, 16456, 16524, 16592, 16660, 16728, 16796, 16864, 16932, 17000, 17068, 17136, 17204, 17272, 17340, 
0, 69, 138, 207, 276, 345, 414, 483, 552, 621, 690, 759, 828, 897, 966, 1035, 1104, 1173, 1242, 1311, 1380, 1449, 1518, 1587, 1656, 1725, 1794, 1863, 1932, 2001, 2070, 2139, 2208, 2277, 2346, 2415, 2484, 2553, 2622, 2691, 2760, 2829, 2898, 2967, 3036, 3105, 3174, 3243, 3312, 3381, 3450, 3519, 3588, 3657, 3726, 3795, 3864, 3933, 4002, 4071, 4140, 4209, 4278, 4347, 4416, 4485, 4554, 4623, 4692, 4761, 4830, 4899, 4968, 5037, 5106, 5175, 5244, 5313, 5382, 5451, 5520, 5589, 5658, 5727, 5796, 5865, 5934, 6003, 6072, 6141, 6210, 6279, 6348, 6417, 6486, 6555, 6624, 6693, 6762, 6831, 6900, 6969, 7038, 7107, 7176, 7245, 7314, 7383, 7452, 7521, 7590, 7659, 7728, 7797, 7866, 7935, 8004, 8073, 8142, 8211, 8280, 8349, 8418, 8487, 8556, 8625, 8694, 8763, 8832, 8901, 8970, 9039, 9108, 9177, 9246, 9315, 9384, 9453, 9522, 9591, 9660, 9729, 9798, 9867, 9936, 10005, 10074, 10143, 10212, 10281, 10350, 10419, 10488, 10557, 10626, 10695, 10764, 10833, 10902, 10971, 11040, 11109, 11178, 11247, 11316, 11385, 11454, 11523, 11592, 11661, 11730, 11799, 11868, 11937, 12006, 12075, 12144, 12213, 12282, 12351, 12420, 12489, 12558, 12627, 12696, 12765, 12834, 12903, 12972, 13041, 13110, 13179, 13248, 13317, 13386, 13455, 13524, 13593, 13662, 13731, 13800, 13869, 13938, 14007, 14076, 14145, 14214, 14283, 14352, 14421, 14490, 14559, 14628, 14697, 14766, 14835, 14904, 14973, 15042, 15111, 15180, 15249, 15318, 15387, 15456, 15525, 15594, 15663, 15732, 15801, 15870, 15939, 16008, 16077, 16146, 16215, 16284, 16353, 16422, 16491, 16560, 16629, 16698, 16767, 16836, 16905, 16974, 17043, 17112, 17181, 17250, 17319, 17388, 17457, 17526, 17595, 
0, 70, 140, 210, 280, 350, 420, 490, 560, 630, 700, 770, 840, 910, 980, 1050, 1120, 1190, 1260, 1330, 1400, 1470, 1540, 1610, 1680, 1750, 1820, 1890, 1960, 2030, 2100, 2170, 2240, 2310, 2380, 2450, 2520, 2590, 2660, 2730, 2800, 2870, 2940, 3010, 3080, 3150, 3220, 3290, 3360, 3430, 3500, 3570, 3640, 3710, 3780, 3850, 3920, 3990, 4060, 4130, 4200, 4270, 4340, 4410, 4480, 4550, 4620, 4690, 4760, 4830, 4900, 4970, 5040, 5110, 5180, 5250, 5320, 5390, 5460, 5530, 5600, 5670, 5740, 5810, 5880, 5950, 6020, 6090, 6160, 6230, 6300, 6370, 6440, 6510, 6580, 6650, 6720, 6790, 6860, 6930, 7000, 7070, 7140, 7210, 7280, 7350, 7420, 7490, 7560, 7630, 7700, 7770, 7840, 7910, 7980, 8050, 8120, 8190, 8260, 8330, 8400, 8470, 8540, 8610, 8680, 8750, 8820, 8890, 8960, 9030, 9100, 9170, 9240, 9310, 9380, 9450, 9520, 9590, 9660, 9730, 9800, 9870, 9940, 10010, 10080, 10150, 10220, 10290, 10360, 10430, 10500, 10570, 10640, 10710, 10780, 10850, 10920, 10990, 11060, 11130, 11200, 11270, 11340, 11410, 11480, 11550, 11620, 11690, 11760, 11830, 11900, 11970, 12040, 12110, 12180, 12250, 12320, 12390, 12460, 12530, 12600, 12670, 12740, 12810, 12880, 12950, 13020, 13090, 13160, 13230, 13300, 13370, 13440, 13510, 13580, 13650, 13720, 13790, 13860, 13930, 14000, 14070, 14140, 14210, 14280, 14350, 14420, 14490, 14560, 14630, 14700, 14770, 14840, 14910, 14980, 15050, 15120, 15190, 15260, 15330, 15400, 15470, 15540, 15610, 15680, 15750, 15820, 15890, 15960, 16030, 16100, 16170, 16240, 16310, 16380, 16450, 16520, 16590, 16660, 16730, 16800, 16870, 16940, 17010, 17080, 17150, 17220, 17290, 17360, 17430, 17500, 17570, 17640, 17710, 17780, 17850, 
0, 71, 142, 213, 284, 355, 426, 497, 568, 639, 710, 781, 852, 923, 994, 1065, 1136, 1207, 1278, 1349, 1420, 1491, 1562, 1633, 1704, 1775, 1846, 1917, 1988, 2059, 2130, 2201, 2272, 2343, 2414, 2485, 2556, 2627, 2698, 2769, 2840, 2911, 2982, 3053, 3124, 3195, 3266, 3337, 3408, 3479, 3550, 3621, 3692, 3763, 3834, 3905, 3976, 4047, 4118, 4189, 4260, 4331, 4402, 4473, 4544, 4615, 4686, 4757, 4828, 4899, 4970, 5041, 5112, 5183, 5254, 5325, 5396, 5467, 5538, 5609, 5680, 5751, 5822, 5893, 5964, 6035, 6106, 6177, 6248, 6319, 6390, 6461, 6532, 6603, 6674, 6745, 6816, 6887, 6958, 7029, 7100, 7171, 7242, 7313, 7384, 7455, 7526, 7597, 7668, 7739, 7810, 7881, 7952, 8023, 8094, 8165, 8236, 8307, 8378, 8449, 8520, 8591, 8662, 8733, 8804, 8875, 8946, 9017, 9088, 9159, 9230, 9301, 9372, 9443, 9514, 9585, 9656, 9727, 9798, 9869, 9940, 10011, 10082, 10153, 10224, 10295, 10366, 10437, 10508, 10579, 10650, 10721, 10792, 10863, 10934, 11005, 11076, 11147, 11218, 11289, 11360, 11431, 11502, 11573, 11644, 11715, 11786, 11857, 11928, 11999, 12070, 12141, 12212, 12283, 12354, 12425, 12496, 12567, 12638, 12709, 12780, 12851, 12922, 12993, 13064, 13135, 13206, 13277, 13348, 13419, 13490, 13561, 13632, 13703, 13774, 13845, 13916, 13987, 14058, 14129, 14200, 14271, 14342, 14413, 14484, 14555, 14626, 14697, 14768, 14839, 14910, 14981, 15052, 15123, 15194, 15265, 15336, 15407, 15478, 15549, 15620, 15691, 15762, 15833, 15904, 15975, 16046, 16117, 16188, 16259, 16330, 16401, 16472, 16543, 16614, 16685, 16756, 16827, 16898, 16969, 17040, 17111, 17182, 17253, 17324, 17395, 17466, 17537, 17608, 17679, 17750, 17821, 17892, 17963, 18034, 18105, 
0, 72, 144, 216, 288, 360, 432, 504, 576, 648, 720, 792, 864, 936, 1008, 1080, 1152, 1224, 1296, 1368, 1440, 1512, 1584, 1656, 1728, 1800, 1872, 1944, 2016, 2088, 2160, 2232, 2304, 2376, 2448, 2520, 2592, 2664, 2736, 2808, 2880, 2952, 3024, 3096, 3168, 3240, 3312, 3384, 3456, 3528, 3600, 3672, 3744, 3816, 3888, 3960, 4032, 4104, 4176, 4248, 4320, 4392, 4464, 4536, 4608, 4680, 4752, 4824, 4896, 4968, 5040, 5112, 5184, 5256, 5328, 5400, 5472, 5544, 5616, 5688, 5760, 5832, 5904, 5976, 6048, 6120, 6192, 6264, 6336, 6408, 6480, 6552, 6624, 6696, 6768, 6840, 6912, 6984, 7056, 7128, 7200, 7272, 7344, 7416, 7488, 7560, 7632, 7704, 7776, 7848, 7920, 7992, 8064, 8136, 8208, 8280, 8352, 8424, 8496, 8568, 8640, 8712, 8784, 8856, 8928, 9000, 9072, 9144, 9216, 9288, 9360, 9432, 9504, 9576, 9648, 9720, 9792, 9864, 9936, 10008, 10080, 10152, 10224, 10296, 10368, 10440, 10512, 10584, 10656, 10728, 10800, 10872, 10944, 11016, 11088, 11160, 11232, 11304, 11376, 11448, 11520, 11592, 11664, 11736, 11808, 11880, 11952, 12024, 12096, 12168, 12240, 12312, 12384, 12456, 12528, 12600, 12672, 12744, 12816, 12888, 12960, 13032, 13104, 13176, 13248, 13320, 13392, 13464, 13536, 13608, 13680, 13752, 13824, 13896, 13968, 14040, 14112, 14184, 14256, 14328, 14400, 14472, 14544, 14616, 14688, 14760, 14832, 14904, 14976, 15048, 15120, 15192, 15264, 15336, 15408, 15480, 15552, 15624, 15696, 15768, 15840, 15912, 15984, 16056, 16128, 16200, 16272, 16344, 16416, 16488, 16560, 16632, 16704, 16776, 16848, 16920, 16992, 17064, 17136, 17208, 17280, 17352, 17424, 17496, 17568, 17640, 17712, 17784, 17856, 17928, 18000, 18072, 18144, 18216, 18288, 18360, 
0, 73, 146, 219, 292, 365, 438, 511, 584, 657, 730, 803, 876, 949, 1022, 1095, 1168, 1241, 1314, 1387, 1460, 1533, 1606, 1679, 1752, 1825, 1898, 1971, 2044, 2117, 2190, 2263, 2336, 2409, 2482, 2555, 2628, 2701, 2774, 2847, 2920, 2993, 3066, 3139, 3212, 3285, 3358, 3431, 3504, 3577, 3650, 3723, 3796, 3869, 3942, 4015, 4088, 4161, 4234, 4307, 4380, 4453, 4526, 4599, 4672, 4745, 4818, 4891, 4964, 5037, 5110, 5183, 5256, 5329, 5402, 5475, 5548, 5621, 5694, 5767, 5840, 5913, 5986, 6059, 6132, 6205, 6278, 6351, 6424, 6497, 6570, 6643, 6716, 6789, 6862, 6935, 7008, 7081, 7154, 7227, 7300, 7373, 7446, 7519, 7592, 7665, 7738, 7811, 7884, 7957, 8030, 8103, 8176, 8249, 8322, 8395, 8468, 8541, 8614, 8687, 8760, 8833, 8906, 8979, 9052, 9125, 9198, 9271, 9344, 9417, 9490, 9563, 9636, 9709, 9782, 9855, 9928, 10001, 10074, 10147, 10220, 10293, 10366, 10439, 10512, 10585, 10658, 10731, 10804, 10877, 10950, 11023, 11096, 11169, 11242, 11315, 11388, 11461, 11534, 11607, 11680, 11753, 11826, 11899, 11972, 12045, 12118, 12191, 12264, 12337, 12410, 12483, 12556, 12629, 12702, 12775, 12848, 12921, 12994, 13067, 13140, 13213, 13286, 13359, 13432, 13505, 13578, 13651, 13724, 13797, 13870, 13943, 14016, 14089, 14162, 14235, 14308, 14381, 14454, 14527, 14600, 14673, 14746, 14819, 14892, 14965, 15038, 15111, 15184, 15257, 15330, 15403, 15476, 15549, 15622, 15695, 15768, 15841, 15914, 15987, 16060, 16133, 16206, 16279, 16352, 16425, 16498, 16571, 16644, 16717, 16790, 16863, 16936, 17009, 17082, 17155, 17228, 17301, 17374, 17447, 17520, 17593, 17666, 17739, 17812, 17885, 17958, 18031, 18104, 18177, 18250, 18323, 18396, 18469, 18542, 18615, 
0, 74, 148, 222, 296, 370, 444, 518, 592, 666, 740, 814, 888, 962, 1036, 1110, 1184, 1258, 1332, 1406, 1480, 1554, 1628, 1702, 1776, 1850, 1924, 1998, 2072, 2146, 2220, 2294, 2368, 2442, 2516, 2590, 2664, 2738, 2812, 2886, 2960, 3034, 3108, 3182, 3256, 3330, 3404, 3478, 3552, 3626, 3700, 3774, 3848, 3922, 3996, 4070, 4144, 4218, 4292, 4366, 4440, 4514, 4588, 4662, 4736, 4810, 4884, 4958, 5032, 5106, 5180, 5254, 5328, 5402, 5476, 5550, 5624, 5698, 5772, 5846, 5920, 5994, 6068, 6142, 6216, 6290, 6364, 6438, 6512, 6586, 6660, 6734, 6808, 6882, 6956, 7030, 7104, 7178, 7252, 7326, 7400, 7474, 7548, 7622, 7696, 7770, 7844, 7918, 7992, 8066, 8140, 8214, 8288, 8362, 8436, 8510, 8584, 8658, 8732, 8806, 8880, 8954, 9028, 9102, 9176, 9250, 9324, 9398, 9472, 9546, 9620, 9694, 9768, 9842, 9916, 9990, 10064, 10138, 10212, 10286, 10360, 10434, 10508, 10582, 10656, 10730, 10804, 10878, 10952, 11026, 11100, 11174, 11248, 11322, 11396, 11470, 11544, 11618, 11692, 11766, 11840, 11914, 11988, 12062, 12136, 12210, 12284, 12358, 12432, 12506, 12580, 12654, 12728, 12802, 12876, 12950, 13024, 13098, 13172, 13246, 13320, 13394, 13468, 13542, 13616, 13690, 13764, 13838, 13912, 13986, 14060, 14134, 14208, 14282, 14356, 14430, 14504, 14578, 14652, 14726, 14800, 14874, 14948, 15022, 15096, 15170, 15244, 15318, 15392, 15466, 15540, 15614, 15688, 15762, 15836, 15910, 15984, 16058, 16132, 16206, 16280, 16354, 16428, 16502, 16576, 16650, 16724, 16798, 16872, 16946, 17020, 17094, 17168, 17242, 17316, 17390, 17464, 17538, 17612, 17686, 17760, 17834, 17908, 17982, 18056, 18130, 18204, 18278, 18352, 18426, 18500, 18574, 18648, 18722, 18796, 18870, 
0, 75, 150, 225, 300, 375, 450, 525, 600, 675, 750, 825, 900, 975, 1050, 1125, 1200, 1275, 1350, 1425, 1500, 1575, 1650, 1725, 1800, 1875, 1950, 2025, 2100, 2175, 2250, 2325, 2400, 2475, 2550, 2625, 2700, 2775, 2850, 2925, 3000, 3075, 3150, 3225, 3300, 3375, 3450, 3525, 3600, 3675, 3750, 3825, 3900, 3975, 4050, 4125, 4200, 4275, 4350, 4425, 4500, 4575, 4650, 4725, 4800, 4875, 4950, 5025, 5100, 5175, 5250, 5325, 5400, 5475, 5550, 5625, 5700, 5775, 5850, 5925, 6000, 6075, 6150, 6225, 6300, 6375, 6450, 6525, 6600, 6675, 6750, 6825, 6900, 6975, 7050, 7125, 7200, 7275, 7350, 7425, 7500, 7575, 7650, 7725, 7800, 7875, 7950, 8025, 8100, 8175, 8250, 8325, 8400, 8475, 8550, 8625, 8700, 8775, 8850, 8925, 9000, 9075, 9150, 9225, 9300, 9375, 9450, 9525, 9600, 9675, 9750, 9825, 9900, 9975, 10050, 10125, 10200, 10275, 10350, 10425, 10500, 10575, 10650, 10725, 10800, 10875, 10950, 11025, 11100, 11175, 11250, 11325, 11400, 11475, 11550, 11625, 11700, 11775, 11850, 11925, 12000, 12075, 12150, 12225, 12300, 12375, 12450, 12525, 12600, 12675, 12750, 12825, 12900, 12975, 13050, 13125, 13200, 13275, 13350, 13425, 13500, 13575, 13650, 13725, 13800, 13875, 13950, 14025, 14100, 14175, 14250, 14325, 14400, 14475, 14550, 14625, 14700, 14775, 14850, 14925, 15000, 15075, 15150, 15225, 15300, 15375, 15450, 15525, 15600, 15675, 15750, 15825, 15900, 15975, 16050, 16125, 16200, 16275, 16350, 16425, 16500, 16575, 16650, 16725, 16800, 16875, 16950, 17025, 17100, 17175, 17250, 17325, 17400, 17475, 17550, 17625, 17700, 17775, 17850, 17925, 18000, 18075, 18150, 18225, 18300, 18375, 18450, 18525, 18600, 18675, 18750, 18825, 18900, 18975, 19050, 19125, 
0, 76, 152, 228, 304, 380, 456, 532, 608, 684, 760, 836, 912, 988, 1064, 1140, 1216, 1292, 1368, 1444, 1520, 1596, 1672, 1748, 1824, 1900, 1976, 2052, 2128, 2204, 2280, 2356, 2432, 2508, 2584, 2660, 2736, 2812, 2888, 2964, 3040, 3116, 3192, 3268, 3344, 3420, 3496, 3572, 3648, 3724, 3800, 3876, 3952, 4028, 4104, 4180, 4256, 4332, 4408, 4484, 4560, 4636, 4712, 4788, 4864, 4940, 5016, 5092, 5168, 5244, 5320, 5396, 5472, 5548, 5624, 5700, 5776, 5852, 5928, 6004, 6080, 6156, 6232, 6308, 6384, 6460, 6536, 6612, 6688, 6764, 6840, 6916, 6992, 7068, 7144, 7220, 7296, 7372, 7448, 7524, 7600, 7676, 7752, 7828, 7904, 7980, 8056, 8132, 8208, 8284, 8360, 8436, 8512, 8588, 8664, 8740, 8816, 8892, 8968, 9044, 9120, 9196, 9272, 9348, 9424, 9500, 9576, 9652, 9728, 9804, 9880, 9956, 10032, 10108, 10184, 10260, 10336, 10412, 10488, 10564, 10640, 10716, 10792, 10868, 10944, 11020, 11096, 11172, 11248, 11324, 11400, 11476, 11552, 11628, 11704, 11780, 11856, 11932, 12008, 12084, 12160, 12236, 12312, 12388, 12464, 12540, 12616, 12692, 12768, 12844, 12920, 12996, 13072, 13148, 13224, 13300, 13376, 13452, 13528, 13604, 13680, 13756, 13832, 13908, 13984, 14060, 14136, 14212, 14288, 14364, 14440, 14516, 14592, 14668, 14744, 14820, 14896, 14972, 15048, 15124, 15200, 15276, 15352, 15428, 15504, 15580, 15656, 15732, 15808, 15884, 15960, 16036, 16112, 16188, 16264, 16340, 16416, 16492, 16568, 16644, 16720, 16796, 16872, 16948, 17024, 17100, 17176, 17252, 17328, 17404, 17480, 17556, 17632, 17708, 17784, 17860, 17936, 18012, 18088, 18164, 18240, 18316, 18392, 18468, 18544, 18620, 18696, 18772, 18848, 18924, 19000, 19076, 19152, 19228, 19304, 19380, 
0, 77, 154, 231, 308, 385, 462, 539, 616, 693, 770, 847, 924, 1001, 1078, 1155, 1232, 1309, 1386, 1463, 1540, 1617, 1694, 1771, 1848, 1925, 2002, 2079, 2156, 2233, 2310, 2387, 2464, 2541, 2618, 2695, 2772, 2849, 2926, 3003, 3080, 3157, 3234, 3311, 3388, 3465, 3542, 3619, 3696, 3773, 3850, 3927, 4004, 4081, 4158, 4235, 4312, 4389, 4466, 4543, 4620, 4697, 4774, 4851, 4928, 5005, 5082, 5159, 5236, 5313, 5390, 5467, 5544, 5621, 5698, 5775, 5852, 5929, 6006, 6083, 6160, 6237, 6314, 6391, 6468, 6545, 6622, 6699, 6776, 6853, 6930, 7007, 7084, 7161, 7238, 7315, 7392, 7469, 7546, 7623, 7700, 7777, 7854, 7931, 8008, 8085, 8162, 8239, 8316, 8393, 8470, 8547, 8624, 8701, 8778, 8855, 8932, 9009, 9086, 9163, 9240, 9317, 9394, 9471, 9548, 9625, 9702, 9779, 9856, 9933, 10010, 10087, 10164, 10241, 10318, 10395, 10472, 10549, 10626, 10703, 10780, 10857, 10934, 11011, 11088, 11165, 11242, 11319, 11396, 11473, 11550, 11627, 11704, 11781, 11858, 11935, 12012, 12089, 12166, 12243, 12320, 12397, 12474, 12551, 12628, 12705, 12782, 12859, 12936, 13013, 13090, 13167, 13244, 13321, 13398, 13475, 13552, 13629, 13706, 13783, 13860, 13937, 14014, 14091, 14168, 14245, 14322, 14399, 14476, 14553, 14630, 14707, 14784, 14861, 14938, 15015, 15092, 15169, 15246, 15323, 15400, 15477, 15554, 15631, 15708, 15785, 15862, 15939, 16016, 16093, 16170, 16247, 16324, 16401, 16478, 16555, 16632, 16709, 16786, 16863, 16940, 17017, 17094, 17171, 17248, 17325, 17402, 17479, 17556, 17633, 17710, 17787, 17864, 17941, 18018, 18095, 18172, 18249, 18326, 18403, 18480, 18557, 18634, 18711, 18788, 18865, 18942, 19019, 19096, 19173, 19250, 19327, 19404, 19481, 19558, 19635, 
0, 78, 156, 234, 312, 390, 468, 546, 624, 702, 780, 858, 936, 1014, 1092, 1170, 1248, 1326, 1404, 1482, 1560, 1638, 1716, 1794, 1872, 1950, 2028, 2106, 2184, 2262, 2340, 2418, 2496, 2574, 2652, 2730, 2808, 2886, 2964, 3042, 3120, 3198, 3276, 3354, 3432, 3510, 3588, 3666, 3744, 3822, 3900, 3978, 4056, 4134, 4212, 4290, 4368, 4446, 4524, 4602, 4680, 4758, 4836, 4914, 4992, 5070, 5148, 5226, 5304, 5382, 5460, 5538, 5616, 5694, 5772, 5850, 5928, 6006, 6084, 6162, 6240, 6318, 6396, 6474, 6552, 6630, 6708, 6786, 6864, 6942, 7020, 7098, 7176, 7254, 7332, 7410, 7488, 7566, 7644, 7722, 7800, 7878, 7956, 8034, 8112, 8190, 8268, 8346, 8424, 8502, 8580, 8658, 8736, 8814, 8892, 8970, 9048, 9126, 9204, 9282, 9360, 9438, 9516, 9594, 9672, 9750, 9828, 9906, 9984, 10062, 10140, 10218, 10296, 10374, 10452, 10530, 10608, 10686, 10764, 10842, 10920, 10998, 11076, 11154, 11232, 11310, 11388, 11466, 11544, 11622, 11700, 11778, 11856, 11934, 12012, 12090, 12168, 12246, 12324, 12402, 12480, 12558, 12636, 12714, 12792, 12870, 12948, 13026, 13104, 13182, 13260, 13338, 13416, 13494, 13572, 13650, 13728, 13806, 13884, 13962, 14040, 14118, 14196, 14274, 14352, 14430, 14508, 14586, 14664, 14742, 14820, 14898, 14976, 15054, 15132, 15210, 15288, 15366, 15444, 15522, 15600, 15678, 15756, 15834, 15912, 15990, 16068, 16146, 16224, 16302, 16380, 16458, 16536, 16614, 16692, 16770, 16848, 16926, 17004, 17082, 17160, 17238, 17316, 17394, 17472, 17550, 17628, 17706, 17784, 17862, 17940, 18018, 18096, 18174, 18252, 18330, 18408, 18486, 18564, 18642, 18720, 18798, 18876, 18954, 19032, 19110, 19188, 19266, 19344, 19422, 19500, 19578, 19656, 19734, 19812, 19890, 
0, 79, 158, 237, 316, 395, 474, 553, 632, 711, 790, 869, 948, 1027, 1106, 1185, 1264, 1343, 1422, 1501, 1580, 1659, 1738, 1817, 1896, 1975, 2054, 2133, 2212, 2291, 2370, 2449, 2528, 2607, 2686, 2765, 2844, 2923, 3002, 3081, 3160, 3239, 3318, 3397, 3476, 3555, 3634, 3713, 3792, 3871, 3950, 4029, 4108, 4187, 4266, 4345, 4424, 4503, 4582, 4661, 4740, 4819, 4898, 4977, 5056, 5135, 5214, 5293, 5372, 5451, 5530, 5609, 5688, 5767, 5846, 5925, 6004, 6083, 6162, 6241, 6320, 6399, 6478, 6557, 6636, 6715, 6794, 6873, 6952, 7031, 7110, 7189, 7268, 7347, 7426, 7505, 7584, 7663, 7742, 7821, 7900, 7979, 8058, 8137, 8216, 8295, 8374, 8453, 8532, 8611, 8690, 8769, 8848, 8927, 9006, 9085, 9164, 9243, 9322, 9401, 9480, 9559, 9638, 9717, 9796, 9875, 9954, 10033, 10112, 10191, 10270, 10349, 10428, 10507, 10586, 10665, 10744, 10823, 10902, 10981, 11060, 11139, 11218, 11297, 11376, 11455, 11534, 11613, 11692, 11771, 11850, 11929, 12008, 12087, 12166, 12245, 12324, 12403, 12482, 12561, 12640, 12719, 12798, 12877, 12956, 13035, 13114, 13193, 13272, 13351, 13430, 13509, 13588, 13667, 13746, 13825, 13904, 13983, 14062, 14141, 14220, 14299, 14378, 14457, 14536, 14615, 14694, 14773, 14852, 14931, 15010, 15089, 15168, 15247, 15326, 15405, 15484, 15563, 15642, 15721, 15800, 15879, 15958, 16037, 16116, 16195, 16274, 16353, 16432, 16511, 16590, 16669, 16748, 16827, 16906, 16985, 17064, 17143, 17222, 17301, 17380, 17459, 17538, 17617, 17696, 17775, 17854, 17933, 18012, 18091, 18170, 18249, 18328, 18407, 18486, 18565, 18644, 18723, 18802, 18881, 18960, 19039, 19118, 19197, 19276, 19355, 19434, 19513, 19592, 19671, 19750, 19829, 19908, 19987, 20066, 20145, 
0, 80, 160, 240, 320, 400, 480, 560, 640, 720, 800, 880, 960, 1040, 1120, 1200, 1280, 1360, 1440, 1520, 1600, 1680, 1760, 1840, 1920, 2000, 2080, 2160, 2240, 2320, 2400, 2480, 2560, 2640, 2720, 2800, 2880, 2960, 3040, 3120, 3200, 3280, 3360, 3440, 3520, 3600, 3680, 3760, 3840, 3920, 4000, 4080, 4160, 4240, 4320, 4400, 4480, 4560, 4640, 4720, 4800, 4880, 4960, 5040, 5120, 5200, 5280, 5360, 5440, 5520, 5600, 5680, 5760, 5840, 5920, 6000, 6080, 6160, 6240, 6320, 6400, 6480, 6560, 6640, 6720, 6800, 6880, 6960, 7040, 7120, 7200, 7280, 7360, 7440, 7520, 7600, 7680, 7760, 7840, 7920, 8000, 8080, 8160, 8240, 8320, 8400, 8480, 8560, 8640, 8720, 8800, 8880, 8960, 9040, 9120, 9200, 9280, 9360, 9440, 9520, 9600, 9680, 9760, 9840, 9920, 10000, 10080, 10160, 10240, 10320, 10400, 10480, 10560, 10640, 10720, 10800, 10880, 10960, 11040, 11120, 11200, 11280, 11360, 11440, 11520, 11600, 11680, 11760, 11840, 11920, 12000, 12080, 12160, 12240, 12320, 12400, 12480, 12560, 12640, 12720, 12800, 12880, 12960, 13040, 13120, 13200, 13280, 13360, 13440, 13520, 13600, 13680, 13760, 13840, 13920, 14000, 14080, 14160, 14240, 14320, 14400, 14480, 14560, 14640, 14720, 14800, 14880, 14960, 15040, 15120, 15200, 15280, 15360, 15440, 15520, 15600, 15680, 15760, 15840, 15920, 16000, 16080, 16160, 16240, 16320, 16400, 16480, 16560, 16640, 16720, 16800, 16880, 16960, 17040, 17120, 17200, 17280, 17360, 17440, 17520, 17600, 17680, 17760, 17840, 17920, 18000, 18080, 18160, 18240, 18320, 18400, 18480, 18560, 18640, 18720, 18800, 18880, 18960, 19040, 19120, 19200, 19280, 19360, 19440, 19520, 19600, 19680, 19760, 19840, 19920, 20000, 20080, 20160, 20240, 20320, 20400, 
0, 81, 162, 243, 324, 405, 486, 567, 648, 729, 810, 891, 972, 1053, 1134, 1215, 1296, 1377, 1458, 1539, 1620, 1701, 1782, 1863, 1944, 2025, 2106, 2187, 2268, 2349, 2430, 2511, 2592, 2673, 2754, 2835, 2916, 2997, 3078, 3159, 3240, 3321, 3402, 3483, 3564, 3645, 3726, 3807, 3888, 3969, 4050, 4131, 4212, 4293, 4374, 4455, 4536, 4617, 4698, 4779, 4860, 4941, 5022, 5103, 5184, 5265, 5346, 5427, 5508, 5589, 5670, 5751, 5832, 5913, 5994, 6075, 6156, 6237, 6318, 6399, 6480, 6561, 6642, 6723, 6804, 6885, 6966, 7047, 7128, 7209, 7290, 7371, 7452, 7533, 7614, 7695, 7776, 7857, 7938, 8019, 8100, 8181, 8262, 8343, 8424, 8505, 8586, 8667, 8748, 8829, 8910, 8991, 9072, 9153, 9234, 9315, 9396, 9477, 9558, 9639, 9720, 9801, 9882, 9963, 10044, 10125, 10206, 10287, 10368, 10449, 10530, 10611, 10692, 10773, 10854, 10935, 11016, 11097, 11178, 11259, 11340, 11421, 11502, 11583, 11664, 11745, 11826, 11907, 11988, 12069, 12150, 12231, 12312, 12393, 12474, 12555, 12636, 12717, 12798, 12879, 12960, 13041, 13122, 13203, 13284, 13365, 13446, 13527, 13608, 13689, 13770, 13851, 13932, 14013, 14094, 14175, 14256, 14337, 14418, 14499, 14580, 14661, 14742, 14823, 14904, 14985, 15066, 15147, 15228, 15309, 15390, 15471, 15552, 15633, 15714, 15795, 15876, 15957, 16038, 16119, 16200, 16281, 16362, 16443, 16524, 16605, 16686, 16767, 16848, 16929, 17010, 17091, 17172, 17253, 17334, 17415, 17496, 17577, 17658, 17739, 17820, 17901, 17982, 18063, 18144, 18225, 18306, 18387, 18468, 18549, 18630, 18711, 18792, 18873, 18954, 19035, 19116, 19197, 19278, 19359, 19440, 19521, 19602, 19683, 19764, 19845, 19926, 20007, 20088, 20169, 20250, 20331, 20412, 20493, 20574, 20655, 
0, 82, 164, 246, 328, 410, 492, 574, 656, 738, 820, 902, 984, 1066, 1148, 1230, 1312, 1394, 1476, 1558, 1640, 1722, 1804, 1886, 1968, 2050, 2132, 2214, 2296, 2378, 2460, 2542, 2624, 2706, 2788, 2870, 2952, 3034, 3116, 3198, 3280, 3362, 3444, 3526, 3608, 3690, 3772, 3854, 3936, 4018, 4100, 4182, 4264, 4346, 4428, 4510, 4592, 4674, 4756, 4838, 4920, 5002, 5084, 5166, 5248, 5330, 5412, 5494, 5576, 5658, 5740, 5822, 5904, 5986, 6068, 6150, 6232, 6314, 6396, 6478, 6560, 6642, 6724, 6806, 6888, 6970, 7052, 7134, 7216, 7298, 7380, 7462, 7544, 7626, 7708, 7790, 7872, 7954, 8036, 8118, 8200, 8282, 8364, 8446, 8528, 8610, 8692, 8774, 8856, 8938, 9020, 9102, 9184, 9266, 9348, 9430, 9512, 9594, 9676, 9758, 9840, 9922, 10004, 10086, 10168, 10250, 10332, 10414, 10496, 10578, 10660, 10742, 10824, 10906, 10988, 11070, 11152, 11234, 11316, 11398, 11480, 11562, 11644, 11726, 11808, 11890, 11972, 12054, 12136, 12218, 12300, 12382, 12464, 12546, 12628, 12710, 12792, 12874, 12956, 13038, 13120, 13202, 13284, 13366, 13448, 13530, 13612, 13694, 13776, 13858, 13940, 14022, 14104, 14186, 14268, 14350, 14432, 14514, 14596, 14678, 14760, 14842, 14924, 15006, 15088, 15170, 15252, 15334, 15416, 15498, 15580, 15662, 15744, 15826, 15908, 15990, 16072, 16154, 16236, 16318, 16400, 16482, 16564, 16646, 16728, 16810, 16892, 16974, 17056, 17138, 17220, 17302, 17384, 17466, 17548, 17630, 17712, 17794, 17876, 17958, 18040, 18122, 18204, 18286, 18368, 18450, 18532, 18614, 18696, 18778, 18860, 18942, 19024, 19106, 19188, 19270, 19352, 19434, 19516, 19598, 19680, 19762, 19844, 19926, 20008, 20090, 20172, 20254, 20336, 20418, 20500, 20582, 20664, 20746, 20828, 20910, 
0, 83, 166, 249, 332, 415, 498, 581, 664, 747, 830, 913, 996, 1079, 1162, 1245, 1328, 1411, 1494, 1577, 1660, 1743, 1826, 1909, 1992, 2075, 2158, 2241, 2324, 2407, 2490, 2573, 2656, 2739, 2822, 2905, 2988, 3071, 3154, 3237, 3320, 3403, 3486, 3569, 3652, 3735, 3818, 3901, 3984, 4067, 4150, 4233, 4316, 4399, 4482, 4565, 4648, 4731, 4814, 4897, 4980, 5063, 5146, 5229, 5312, 5395, 5478, 5561, 5644, 5727, 5810, 5893, 5976, 6059, 6142, 6225, 6308, 6391, 6474, 6557, 6640, 6723, 6806, 6889, 6972, 7055, 7138, 7221, 7304, 7387, 7470, 7553, 7636, 7719, 7802, 7885, 7968, 8051, 8134, 8217, 8300, 8383, 8466, 8549, 8632, 8715, 8798, 8881, 8964, 9047, 9130, 9213, 9296, 9379, 9462, 9545, 9628, 9711, 9794, 9877, 9960, 10043, 10126, 10209, 10292, 10375, 10458, 10541, 10624, 10707, 10790, 10873, 10956, 11039, 11122, 11205, 11288, 11371, 11454, 11537, 11620, 11703, 11786, 11869, 11952, 12035, 12118, 12201, 12284, 12367, 12450, 12533, 12616, 12699, 12782, 12865, 12948, 13031, 13114, 13197, 13280, 13363, 13446, 13529, 13612, 13695, 13778, 13861, 13944, 14027, 14110, 14193, 14276, 14359, 14442, 14525, 14608, 14691, 14774, 14857, 14940, 15023, 15106, 15189, 15272, 15355, 15438, 15521, 15604, 15687, 15770, 15853, 15936, 16019, 16102, 16185, 16268, 16351, 16434, 16517, 16600, 16683, 16766, 16849, 16932, 17015, 17098, 17181, 17264, 17347, 17430, 17513, 17596, 17679, 17762, 17845, 17928, 18011, 18094, 18177, 18260, 18343, 18426, 18509, 18592, 18675, 18758, 18841, 18924, 19007, 19090, 19173, 19256, 19339, 19422, 19505, 19588, 19671, 19754, 19837, 19920, 20003, 20086, 20169, 20252, 20335, 20418, 20501, 20584, 20667, 20750, 20833, 20916, 20999, 21082, 21165, 
0, 84, 168, 252, 336, 420, 504, 588, 672, 756, 840, 924, 1008, 1092, 1176, 1260, 1344, 1428, 1512, 1596, 1680, 1764, 1848, 1932, 2016, 2100, 2184, 2268, 2352, 2436, 2520, 2604, 2688, 2772, 2856, 2940, 3024, 3108, 3192, 3276, 3360, 3444, 3528, 3612, 3696, 3780, 3864, 3948, 4032, 4116, 4200, 4284, 4368, 4452, 4536, 4620, 4704, 4788, 4872, 4956, 5040, 5124, 5208, 5292, 5376, 5460, 5544, 5628, 5712, 5796, 5880, 5964, 6048, 6132, 6216, 6300, 6384, 6468, 6552, 6636, 6720, 6804, 6888, 6972, 7056, 7140, 7224, 7308, 7392, 7476, 7560, 7644, 7728, 7812, 7896, 7980, 8064, 8148, 8232, 8316, 8400, 8484, 8568, 8652, 8736, 8820, 8904, 8988, 9072, 9156, 9240, 9324, 9408, 9492, 9576, 9660, 9744, 9828, 9912, 9996, 10080, 10164, 10248, 10332, 10416, 10500, 10584, 10668, 10752, 10836, 10920, 11004, 11088, 11172, 11256, 11340, 11424, 11508, 11592, 11676, 11760, 11844, 11928, 12012, 12096, 12180, 12264, 12348, 12432, 12516, 12600, 12684, 12768, 12852, 12936, 13020, 13104, 13188, 13272, 13356, 13440, 13524, 13608, 13692, 13776, 13860, 13944, 14028, 14112, 14196, 14280, 14364, 14448, 14532, 14616, 14700, 14784, 14868, 14952, 15036, 15120, 15204, 15288, 15372, 15456, 15540, 15624, 15708, 15792, 15876, 15960, 16044, 16128, 16212, 16296, 16380, 16464, 16548, 16632, 16716, 16800, 16884, 16968, 17052, 17136, 17220, 17304, 17388, 17472, 17556, 17640, 17724, 17808, 17892, 17976, 18060, 18144, 18228, 18312, 18396, 18480, 18564, 18648, 18732, 18816, 18900, 18984, 19068, 19152, 19236, 19320, 19404, 19488, 19572, 19656, 19740, 19824, 19908, 19992, 20076, 20160, 20244, 20328, 20412, 20496, 20580, 20664, 20748, 20832, 20916, 21000, 21084, 21168, 21252, 21336, 21420, 
0, 85, 170, 255, 340, 425, 510, 595, 680, 765, 850, 935, 1020, 1105, 1190, 1275, 1360, 1445, 1530, 1615, 1700, 1785, 1870, 1955, 2040, 2125, 2210, 2295, 2380, 2465, 2550, 2635, 2720, 2805, 2890, 2975, 3060, 3145, 3230, 3315, 3400, 3485, 3570, 3655, 3740, 3825, 3910, 3995, 4080, 4165, 4250, 4335, 4420, 4505, 4590, 4675, 4760, 4845, 4930, 5015, 5100, 5185, 5270, 5355, 5440, 5525, 5610, 5695, 5780, 5865, 5950, 6035, 6120, 6205, 6290, 6375, 6460, 6545, 6630, 6715, 6800, 6885, 6970, 7055, 7140, 7225, 7310, 7395, 7480, 7565, 7650, 7735, 7820, 7905, 7990, 8075, 8160, 8245, 8330, 8415, 8500, 8585, 8670, 8755, 8840, 8925, 9010, 9095, 9180, 9265, 9350, 9435, 9520, 9605, 9690, 9775, 9860, 9945, 10030, 10115, 10200, 10285, 10370, 10455, 10540, 10625, 10710, 10795, 10880, 10965, 11050, 11135, 11220, 11305, 11390, 11475, 11560, 11645, 11730, 11815, 11900, 11985, 12070, 12155, 12240, 12325, 12410, 12495, 12580, 12665, 12750, 12835, 12920, 13005, 13090, 13175, 13260, 13345, 13430, 13515, 13600, 13685, 13770, 13855, 13940, 14025, 14110, 14195, 14280, 14365, 14450, 14535, 14620, 14705, 14790, 14875, 14960, 15045, 15130, 15215, 15300, 15385, 15470, 15555, 15640, 15725, 15810, 15895, 15980, 16065, 16150, 16235, 16320, 16405, 16490, 16575, 16660, 16745, 16830, 16915, 17000, 17085, 17170, 17255, 17340, 17425, 17510, 17595, 17680, 17765, 17850, 17935, 18020, 18105, 18190, 18275, 18360, 18445, 18530, 18615, 18700, 18785, 18870, 18955, 19040, 19125, 19210, 19295, 19380, 19465, 19550, 19635, 19720, 19805, 19890, 19975, 20060, 20145, 20230, 20315, 20400, 20485, 20570, 20655, 20740, 20825, 20910, 20995, 21080, 21165, 21250, 21335, 21420, 21505, 21590, 21675, 
0, 86, 172, 258, 344, 430, 516, 602, 688, 774, 860, 946, 1032, 1118, 1204, 1290, 1376, 1462, 1548, 1634, 1720, 1806, 1892, 1978, 2064, 2150, 2236, 2322, 2408, 2494, 2580, 2666, 2752, 2838, 2924, 3010, 3096, 3182, 3268, 3354, 3440, 3526, 3612, 3698, 3784, 3870, 3956, 4042, 4128, 4214, 4300, 4386, 4472, 4558, 4644, 4730, 4816, 4902, 4988, 5074, 5160, 5246, 5332, 5418, 5504, 5590, 5676, 5762, 5848, 5934, 6020, 6106, 6192, 6278, 6364, 6450, 6536, 6622, 6708, 6794, 6880, 6966, 7052, 7138, 7224, 7310, 7396, 7482, 7568, 7654, 7740, 7826, 7912, 7998, 8084, 8170, 8256, 8342, 8428, 8514, 8600, 8686, 8772, 8858, 8944, 9030, 9116, 9202, 9288, 9374, 9460, 9546, 9632, 9718, 9804, 9890, 9976, 10062, 10148, 10234, 10320, 10406, 10492, 10578, 10664, 10750, 10836, 10922, 11008, 11094, 11180, 11266, 11352, 11438, 11524, 11610, 11696, 11782, 11868, 11954, 12040, 12126, 12212, 12298, 12384, 12470, 12556, 12642, 12728, 12814, 12900, 12986, 13072, 13158, 13244, 13330, 13416, 13502, 13588, 13674, 13760, 13846, 13932, 14018, 14104, 14190, 14276, 14362, 14448, 14534, 14620, 14706, 14792, 14878, 14964, 15050, 15136, 15222, 15308, 15394, 15480, 15566, 15652, 15738, 15824, 15910, 15996, 16082, 16168, 16254, 16340, 16426, 16512, 16598, 16684, 16770, 16856, 16942, 17028, 17114, 17200, 17286, 17372, 17458, 17544, 17630, 17716, 17802, 17888, 17974, 18060, 18146, 18232, 18318, 18404, 18490, 18576, 18662, 18748, 18834, 18920, 19006, 19092, 19178, 19264, 19350, 19436, 19522, 19608, 19694, 19780, 19866, 19952, 20038, 20124, 20210, 20296, 20382, 20468, 20554, 20640, 20726, 20812, 20898, 20984, 21070, 21156, 21242, 21328, 21414, 21500, 21586, 21672, 21758, 21844, 21930, 
0, 87, 174, 261, 348, 435, 522, 609, 696, 783, 870, 957, 1044, 1131, 1218, 1305, 1392, 1479, 1566, 1653, 1740, 1827, 1914, 2001, 2088, 2175, 2262, 2349, 2436, 2523, 2610, 2697, 2784, 2871, 2958, 3045, 3132, 3219, 3306, 3393, 3480, 3567, 3654, 3741, 3828, 3915, 4002, 4089, 4176, 4263, 4350, 4437, 4524, 4611, 4698, 4785, 4872, 4959, 5046, 5133, 5220, 5307, 5394, 5481, 5568, 5655, 5742, 5829, 5916, 6003, 6090, 6177, 6264, 6351, 6438, 6525, 6612, 6699, 6786, 6873, 6960, 7047, 7134, 7221, 7308, 7395, 7482, 7569, 7656, 7743, 7830, 7917, 8004, 8091, 8178, 8265, 8352, 8439, 8526, 8613, 8700, 8787, 8874, 8961, 9048, 9135, 9222, 9309, 9396, 9483, 9570, 9657, 9744, 9831, 9918, 10005, 10092, 10179, 10266, 10353, 10440, 10527, 10614, 10701, 10788, 10875, 10962, 11049, 11136, 11223, 11310, 11397, 11484, 11571, 11658, 11745, 11832, 11919, 12006, 12093, 12180, 12267, 12354, 12441, 12528, 12615, 12702, 12789, 12876, 12963, 13050, 13137, 13224, 13311, 13398, 13485, 13572, 13659, 13746, 13833, 13920, 14007, 14094, 14181, 14268, 14355, 14442, 14529, 14616, 14703, 14790, 14877, 14964, 15051, 15138, 15225, 15312, 15399, 15486, 15573, 15660, 15747, 15834, 15921, 16008, 16095, 16182, 16269, 16356, 16443, 16530, 16617, 16704, 16791, 16878, 16965, 17052, 17139, 17226, 17313, 17400, 17487, 17574, 17661, 17748, 17835, 17922, 18009, 18096, 18183, 18270, 18357, 18444, 18531, 18618, 18705, 18792, 18879, 18966, 19053, 19140, 19227, 19314, 19401, 19488, 19575, 19662, 19749, 19836, 19923, 20010, 20097, 20184, 20271, 20358, 20445, 20532, 20619, 20706, 20793, 20880, 20967, 21054, 21141, 21228, 21315, 21402, 21489, 21576, 21663, 21750, 21837, 21924, 22011, 22098, 22185, 
0, 88, 176, 264, 352, 440, 528, 616, 704, 792, 880, 968, 1056, 1144, 1232, 1320, 1408, 1496, 1584, 1672, 1760, 1848, 1936, 2024, 2112, 2200, 2288, 2376, 2464, 2552, 2640, 2728, 2816, 2904, 2992, 3080, 3168, 3256, 3344, 3432, 3520, 3608, 3696, 3784, 3872, 3960, 4048, 4136, 4224, 4312, 4400, 4488, 4576, 4664, 4752, 4840, 4928, 5016, 5104, 5192, 5280, 5368, 5456, 5544, 5632, 5720, 5808, 5896, 5984, 6072, 6160, 6248, 6336, 6424, 6512, 6600, 6688, 6776, 6864, 6952, 7040, 7128, 7216, 7304, 7392, 7480, 7568, 7656, 7744, 7832, 7920, 8008, 8096, 8184, 8272, 8360, 8448, 8536, 8624, 8712, 8800, 8888, 8976, 9064, 9152, 9240, 9328, 9416, 9504, 9592, 9680, 9768, 9856, 9944, 10032, 10120, 10208, 10296, 10384, 10472, 10560, 10648, 10736, 10824, 10912, 11000, 11088, 11176, 11264, 11352, 11440, 11528, 11616, 11704, 11792, 11880, 11968, 12056, 12144, 12232, 12320, 12408, 12496, 12584, 12672, 12760, 12848, 12936, 13024, 13112, 13200, 13288, 13376, 13464, 13552, 13640, 13728, 13816, 13904, 13992, 14080, 14168, 14256, 14344, 14432, 14520, 14608, 14696, 14784, 14872, 14960, 15048, 15136, 15224, 15312, 15400, 15488, 15576, 15664, 15752, 15840, 15928, 16016, 16104, 16192, 16280, 16368, 16456, 16544, 16632, 16720, 16808, 16896, 16984, 17072, 17160, 17248, 17336, 17424, 17512, 17600, 17688, 17776, 17864, 17952, 18040, 18128, 18216, 18304, 18392, 18480, 18568, 18656, 18744, 18832, 18920, 19008, 19096, 19184, 19272, 19360, 19448, 19536, 19624, 19712, 19800, 19888, 19976, 20064, 20152, 20240, 20328, 20416, 20504, 20592, 20680, 20768, 20856, 20944, 21032, 21120, 21208, 21296, 21384, 21472, 21560, 21648, 21736, 21824, 21912, 22000, 22088, 22176, 22264, 22352, 22440, 
0, 89, 178, 267, 356, 445, 534, 623, 712, 801, 890, 979, 1068, 1157, 1246, 1335, 1424, 1513, 1602, 1691, 1780, 1869, 1958, 2047, 2136, 2225, 2314, 2403, 2492, 2581, 2670, 2759, 2848, 2937, 3026, 3115, 3204, 3293, 3382, 3471, 3560, 3649, 3738, 3827, 3916, 4005, 4094, 4183, 4272, 4361, 4450, 4539, 4628, 4717, 4806, 4895, 4984, 5073, 5162, 5251, 5340, 5429, 5518, 5607, 5696, 5785, 5874, 5963, 6052, 6141, 6230, 6319, 6408, 6497, 6586, 6675, 6764, 6853, 6942, 7031, 7120, 7209, 7298, 7387, 7476, 7565, 7654, 7743, 7832, 7921, 8010, 8099, 8188, 8277, 8366, 8455, 8544, 8633, 8722, 8811, 8900, 8989, 9078, 9167, 9256, 9345, 9434, 9523, 9612, 9701, 9790, 9879, 9968, 10057, 10146, 10235, 10324, 10413, 10502, 10591, 10680, 10769, 10858, 10947, 11036, 11125, 11214, 11303, 11392, 11481, 11570, 11659, 11748, 11837, 11926, 12015, 12104, 12193, 12282, 12371, 12460, 12549, 12638, 12727, 12816, 12905, 12994, 13083, 13172, 13261, 13350, 13439, 13528, 13617, 13706, 13795, 13884, 13973, 14062, 14151, 14240, 14329, 14418, 14507, 14596, 14685, 14774, 14863, 14952, 15041, 15130, 15219, 15308, 15397, 15486, 15575, 15664, 15753, 15842, 15931, 16020, 16109, 16198, 16287, 16376, 16465, 16554, 16643, 16732, 16821, 16910, 16999, 17088, 17177, 17266, 17355, 17444, 17533, 17622, 17711, 17800, 17889, 17978, 18067, 18156, 18245, 18334, 18423, 18512, 18601, 18690, 18779, 18868, 18957, 19046, 19135, 19224, 19313, 19402, 19491, 19580, 19669, 19758, 19847, 19936, 20025, 20114, 20203, 20292, 20381, 20470, 20559, 20648, 20737, 20826, 20915, 21004, 21093, 21182, 21271, 21360, 21449, 21538, 21627, 21716, 21805, 21894, 21983, 22072, 22161, 22250, 22339, 22428, 22517, 22606, 22695, 
0, 90, 180, 270, 360, 450, 540, 630, 720, 810, 900, 990, 1080, 1170, 1260, 1350, 1440, 1530, 1620, 1710, 1800, 1890, 1980, 2070, 2160, 2250, 2340, 2430, 2520, 2610, 2700, 2790, 2880, 2970, 3060, 3150, 3240, 3330, 3420, 3510, 3600, 3690, 3780, 3870, 3960, 4050, 4140, 4230, 4320, 4410, 4500, 4590, 4680, 4770, 4860, 4950, 5040, 5130, 5220, 5310, 5400, 5490, 5580, 5670, 5760, 5850, 5940, 6030, 6120, 6210, 6300, 6390, 6480, 6570, 6660, 6750, 6840, 6930, 7020, 7110, 7200, 7290, 7380, 7470, 7560, 7650, 7740, 7830, 7920, 8010, 8100, 8190, 8280, 8370, 8460, 8550, 8640, 8730, 8820, 8910, 9000, 9090, 9180, 9270, 9360, 9450, 9540, 9630, 9720, 9810, 9900, 9990, 10080, 10170, 10260, 10350, 10440, 10530, 10620, 10710, 10800, 10890, 10980, 11070, 11160, 11250, 11340, 11430, 11520, 11610, 11700, 11790, 11880, 11970, 12060, 12150, 12240, 12330, 12420, 12510, 12600, 12690, 12780, 12870, 12960, 13050, 13140, 13230, 13320, 13410, 13500, 13590, 13680, 13770, 13860, 13950, 14040, 14130, 14220, 14310, 14400, 14490, 14580, 14670, 14760, 14850, 14940, 15030, 15120, 15210, 15300, 15390, 15480, 15570, 15660, 15750, 15840, 15930, 16020, 16110, 16200, 16290, 16380, 16470, 16560, 16650, 16740, 16830, 16920, 17010, 17100, 17190, 17280, 17370, 17460, 17550, 17640, 17730, 17820, 17910, 18000, 18090, 18180, 18270, 18360, 18450, 18540, 18630, 18720, 18810, 18900, 18990, 19080, 19170, 19260, 19350, 19440, 19530, 19620, 19710, 19800, 19890, 19980, 20070, 20160, 20250, 20340, 20430, 20520, 20610, 20700, 20790, 20880, 20970, 21060, 21150, 21240, 21330, 21420, 21510, 21600, 21690, 21780, 21870, 21960, 22050, 22140, 22230, 22320, 22410, 22500, 22590, 22680, 22770, 22860, 22950, 
0, 91, 182, 273, 364, 455, 546, 637, 728, 819, 910, 1001, 1092, 1183, 1274, 1365, 1456, 1547, 1638, 1729, 1820, 1911, 2002, 2093, 2184, 2275, 2366, 2457, 2548, 2639, 2730, 2821, 2912, 3003, 3094, 3185, 3276, 3367, 3458, 3549, 3640, 3731, 3822, 3913, 4004, 4095, 4186, 4277, 4368, 4459, 4550, 4641, 4732, 4823, 4914, 5005, 5096, 5187, 5278, 5369, 5460, 5551, 5642, 5733, 5824, 5915, 6006, 6097, 6188, 6279, 6370, 6461, 6552, 6643, 6734, 6825, 6916, 7007, 7098, 7189, 7280, 7371, 7462, 7553, 7644, 7735, 7826, 7917, 8008, 8099, 8190, 8281, 8372, 8463, 8554, 8645, 8736, 8827, 8918, 9009, 9100, 9191, 9282, 9373, 9464, 9555, 9646, 9737, 9828, 9919, 10010, 10101, 10192, 10283, 10374, 10465, 10556, 10647, 10738, 10829, 10920, 11011, 11102, 11193, 11284, 11375, 11466, 11557, 11648, 11739, 11830, 11921, 12012, 12103, 12194, 12285, 12376, 12467, 12558, 12649, 12740, 12831, 12922, 13013, 13104, 13195, 13286, 13377, 13468, 13559, 13650, 13741, 13832, 13923, 14014, 14105, 14196, 14287, 14378, 14469, 14560, 14651, 14742, 14833, 14924, 15015, 15106, 15197, 15288, 15379, 15470, 15561, 15652, 15743, 15834, 15925, 16016, 16107, 16198, 16289, 16380, 16471, 16562, 16653, 16744, 16835, 16926, 17017, 17108, 17199, 17290, 17381, 17472, 17563, 17654, 17745, 17836, 17927, 18018, 18109, 18200, 18291, 18382, 18473, 18564, 18655, 18746, 18837, 18928, 19019, 19110, 19201, 19292, 19383, 19474, 19565, 19656, 19747, 19838, 19929, 20020, 20111, 20202, 20293, 20384, 20475, 20566, 20657, 20748, 20839, 20930, 21021, 21112, 21203, 21294, 21385, 21476, 21567, 21658, 21749, 21840, 21931, 22022, 22113, 22204, 22295, 22386, 22477, 22568, 22659, 22750, 22841, 22932, 23023, 23114, 23205, 
0, 92, 184, 276, 368, 460, 552, 644, 736, 828, 920, 1012, 1104, 1196, 1288, 1380, 1472, 1564, 1656, 1748, 1840, 1932, 2024, 2116, 2208, 2300, 2392, 2484, 2576, 2668, 2760, 2852, 2944, 3036, 3128, 3220, 3312, 3404, 3496, 3588, 3680, 3772, 3864, 3956, 4048, 4140, 4232, 4324, 4416, 4508, 4600, 4692, 4784, 4876, 4968, 5060, 5152, 5244, 5336, 5428, 5520, 5612, 5704, 5796, 5888, 5980, 6072, 6164, 6256, 6348, 6440, 6532, 6624, 6716, 6808, 6900, 6992, 7084, 7176, 7268, 7360, 7452, 7544, 7636, 7728, 7820, 7912, 8004, 8096, 8188, 8280, 8372, 8464, 8556, 8648, 8740, 8832, 8924, 9016, 9108, 9200, 9292, 9384, 9476, 9568, 9660, 9752, 9844, 9936, 10028, 10120, 10212, 10304, 10396, 10488, 10580, 10672, 10764, 10856, 10948, 11040, 11132, 11224, 11316, 11408, 11500, 11592, 11684, 11776, 11868, 11960, 12052, 12144, 12236, 12328, 12420, 12512, 12604, 12696, 12788, 12880, 12972, 13064, 13156, 13248, 13340, 13432, 13524, 13616, 13708, 13800, 13892, 13984, 14076, 14168, 14260, 14352, 14444, 14536, 14628, 14720, 14812, 14904, 14996, 15088, 15180, 15272, 15364, 15456, 15548, 15640, 15732, 15824, 15916, 16008, 16100, 16192, 16284, 16376, 16468, 16560, 16652, 16744, 16836, 16928, 17020, 17112, 17204, 17296, 17388, 17480, 17572, 17664, 17756, 17848, 17940, 18032, 18124, 18216, 18308, 18400, 18492, 18584, 18676, 18768, 18860, 18952, 19044, 19136, 19228, 19320, 19412, 19504, 19596, 19688, 19780, 19872, 19964, 20056, 20148, 20240, 20332, 20424, 20516, 20608, 20700, 20792, 20884, 20976, 21068, 21160, 21252, 21344, 21436, 21528, 21620, 21712, 21804, 21896, 21988, 22080, 22172, 22264, 22356, 22448, 22540, 22632, 22724, 22816, 22908, 23000, 23092, 23184, 23276, 23368, 23460, 
0, 93, 186, 279, 372, 465, 558, 651, 744, 837, 930, 1023, 1116, 1209, 1302, 1395, 1488, 1581, 1674, 1767, 1860, 1953, 2046, 2139, 2232, 2325, 2418, 2511, 2604, 2697, 2790, 2883, 2976, 3069, 3162, 3255, 3348, 3441, 3534, 3627, 3720, 3813, 3906, 3999, 4092, 4185, 4278, 4371, 4464, 4557, 4650, 4743, 4836, 4929, 5022, 5115, 5208, 5301, 5394, 5487, 5580, 5673, 5766, 5859, 5952, 6045, 6138, 6231, 6324, 6417, 6510, 6603, 6696, 6789, 6882, 6975, 7068, 7161, 7254, 7347, 7440, 7533, 7626, 7719, 7812, 7905, 7998, 8091, 8184, 8277, 8370, 8463, 8556, 8649, 8742, 8835, 8928, 9021, 9114, 9207, 9300, 9393, 9486, 9579, 9672, 9765, 9858, 9951, 10044, 10137, 10230, 10323, 10416, 10509, 10602, 10695, 10788, 10881, 10974, 11067, 11160, 11253, 11346, 11439, 11532, 11625, 11718, 11811, 11904, 11997, 12090, 12183, 12276, 12369, 12462, 12555, 12648, 12741, 12834, 12927, 13020, 13113, 13206, 13299, 13392, 13485, 13578, 13671, 13764, 13857, 13950, 14043, 14136, 14229, 14322, 14415, 14508, 14601, 14694, 14787, 14880, 14973, 15066, 15159, 15252, 15345, 15438, 15531, 15624, 15717, 15810, 15903, 15996, 16089, 16182, 16275, 16368, 16461, 16554, 16647, 16740, 16833, 16926, 17019, 17112, 17205, 17298, 17391, 17484, 17577, 17670, 17763, 17856, 17949, 18042, 18135, 18228, 18321, 18414, 18507, 18600, 18693, 18786, 18879, 18972, 19065, 19158, 19251, 19344, 19437, 19530, 19623, 19716, 19809, 19902, 19995, 20088, 20181, 20274, 20367, 20460, 20553, 20646, 20739, 20832, 20925, 21018, 21111, 21204, 21297, 21390, 21483, 21576, 21669, 21762, 21855, 21948, 22041, 22134, 22227, 22320, 22413, 22506, 22599, 22692, 22785, 22878, 22971, 23064, 23157, 23250, 23343, 23436, 23529, 23622, 23715, 
0, 94, 188, 282, 376, 470, 564, 658, 752, 846, 940, 1034, 1128, 1222, 1316, 1410, 1504, 1598, 1692, 1786, 1880, 1974, 2068, 2162, 2256, 2350, 2444, 2538, 2632, 2726, 2820, 2914, 3008, 3102, 3196, 3290, 3384, 3478, 3572, 3666, 3760, 3854, 3948, 4042, 4136, 4230, 4324, 4418, 4512, 4606, 4700, 4794, 4888, 4982, 5076, 5170, 5264, 5358, 5452, 5546, 5640, 5734, 5828, 5922, 6016, 6110, 6204, 6298, 6392, 6486, 6580, 6674, 6768, 6862, 6956, 7050, 7144, 7238, 7332, 7426, 7520, 7614, 7708, 7802, 7896, 7990, 8084, 8178, 8272, 8366, 8460, 8554, 8648, 8742, 8836, 8930, 9024, 9118, 9212, 9306, 9400, 9494, 9588, 9682, 9776, 9870, 9964, 10058, 10152, 10246, 10340, 10434, 10528, 10622, 10716, 10810, 10904, 10998, 11092, 11186, 11280, 11374, 11468, 11562, 11656, 11750, 11844, 11938, 12032, 12126, 12220, 12314, 12408, 12502, 12596, 12690, 12784, 12878, 12972, 13066, 13160, 13254, 13348, 13442, 13536, 13630, 13724, 13818, 13912, 14006, 14100, 14194, 14288, 14382, 14476, 14570, 14664, 14758, 14852, 14946, 15040, 15134, 15228, 15322, 15416, 15510, 15604, 15698, 15792, 15886, 15980, 16074, 16168, 16262, 16356, 16450, 16544, 16638, 16732, 16826, 16920, 17014, 17108, 17202, 17296, 17390, 17484, 17578, 17672, 17766, 17860, 17954, 18048, 18142, 18236, 18330, 18424, 18518, 18612, 18706, 18800, 18894, 18988, 19082, 19176, 19270, 19364, 19458, 19552, 19646, 19740, 19834, 19928, 20022, 20116, 20210, 20304, 20398, 20492, 20586, 20680, 20774, 20868, 20962, 21056, 21150, 21244, 21338, 21432, 21526, 21620, 21714, 21808, 21902, 21996, 22090, 22184, 22278, 22372, 22466, 22560, 22654, 22748, 22842, 22936, 23030, 23124, 23218, 23312, 23406, 23500, 23594, 23688, 23782, 23876, 23970, 
0, 95, 190, 285, 380, 475, 570, 665, 760, 855, 950, 1045, 1140, 1235, 1330, 1425, 1520, 1615, 1710, 1805, 1900, 1995, 2090, 2185, 2280, 2375, 2470, 2565, 2660, 2755, 2850, 2945, 3040, 3135, 3230, 3325, 3420, 3515, 3610, 3705, 3800, 3895, 3990, 4085, 4180, 4275, 4370, 4465, 4560, 4655, 4750, 4845, 4940, 5035, 5130, 5225, 5320, 5415, 5510, 5605, 5700, 5795, 5890, 5985, 6080, 6175, 6270, 6365, 6460, 6555, 6650, 6745, 6840, 6935, 7030, 7125, 7220, 7315, 7410, 7505, 7600, 7695, 7790, 7885, 7980, 8075, 8170, 8265, 8360, 8455, 8550, 8645, 8740, 8835, 8930, 9025, 9120, 9215, 9310, 9405, 9500, 9595, 9690, 9785, 9880, 9975, 10070, 10165, 10260, 10355, 10450, 10545, 10640, 10735, 10830, 10925, 11020, 11115, 11210, 11305, 11400, 11495, 11590, 11685, 11780, 11875, 11970, 12065, 12160, 12255, 12350, 12445, 12540, 12635, 12730, 12825, 12920, 13015, 13110, 13205, 13300, 13395, 13490, 13585, 13680, 13775, 13870, 13965, 14060, 14155, 14250, 14345, 14440, 14535, 14630, 14725, 14820, 14915, 15010, 15105, 15200, 15295, 15390, 15485, 15580, 15675, 15770, 15865, 15960, 16055, 16150, 16245, 16340, 16435, 16530, 16625, 16720, 16815, 16910, 17005, 17100, 17195, 17290, 17385, 17480, 17575, 17670, 17765, 17860, 17955, 18050, 18145, 18240, 18335, 18430, 18525, 18620, 18715, 18810, 18905, 19000, 19095, 19190, 19285, 19380, 19475, 19570, 19665, 19760, 19855, 19950, 20045, 20140, 20235, 20330, 20425, 20520, 20615, 20710, 20805, 20900, 20995, 21090, 21185, 21280, 21375, 21470, 21565, 21660, 21755, 21850, 21945, 22040, 22135, 22230, 22325, 22420, 22515, 22610, 22705, 22800, 22895, 22990, 23085, 23180, 23275, 23370, 23465, 23560, 23655, 23750, 23845, 23940, 24035, 24130, 24225, 
0, 96, 192, 288, 384, 480, 576, 672, 768, 864, 960, 1056, 1152, 1248, 1344, 1440, 1536, 1632, 1728, 1824, 1920, 2016, 2112, 2208, 2304, 2400, 2496, 2592, 2688, 2784, 2880, 2976, 3072, 3168, 3264, 3360, 3456, 3552, 3648, 3744, 3840, 3936, 4032, 4128, 4224, 4320, 4416, 4512, 4608, 4704, 4800, 4896, 4992, 5088, 5184, 5280, 5376, 5472, 5568, 5664, 5760, 5856, 5952, 6048, 6144, 6240, 6336, 6432, 6528, 6624, 6720, 6816, 6912, 7008, 7104, 7200, 7296, 7392, 7488, 7584, 7680, 7776, 7872, 7968, 8064, 8160, 8256, 8352, 8448, 8544, 8640, 8736, 8832, 8928, 9024, 9120, 9216, 9312, 9408, 9504, 9600, 9696, 9792, 9888, 9984, 10080, 10176, 10272, 10368, 10464, 10560, 10656, 10752, 10848, 10944, 11040, 11136, 11232, 11328, 11424, 11520, 11616, 11712, 11808, 11904, 12000, 12096, 12192, 12288, 12384, 12480, 12576, 12672, 12768, 12864, 12960, 13056, 13152, 13248, 13344, 13440, 13536, 13632, 13728, 13824, 13920, 14016, 14112, 14208, 14304, 14400, 14496, 14592, 14688, 14784, 14880, 14976, 15072, 15168, 15264, 15360, 15456, 15552, 15648, 15744, 15840, 15936, 16032, 16128, 16224, 16320, 16416, 16512, 16608, 16704, 16800, 16896, 16992, 17088, 17184, 17280, 17376, 17472, 17568, 17664, 17760, 17856, 17952, 18048, 18144, 18240, 18336, 18432, 18528, 18624, 18720, 18816, 18912, 19008, 19104, 19200, 19296, 19392, 19488, 19584, 19680, 19776, 19872, 19968, 20064, 20160, 20256, 20352, 20448, 20544, 20640, 20736, 20832, 20928, 21024, 21120, 21216, 21312, 21408, 21504, 21600, 21696, 21792, 21888, 21984, 22080, 22176, 22272, 22368, 22464, 22560, 22656, 22752, 22848, 22944, 23040, 23136, 23232, 23328, 23424, 23520, 23616, 23712, 23808, 23904, 24000, 24096, 24192, 24288, 24384, 24480, 
0, 97, 194, 291, 388, 485, 582, 679, 776, 873, 970, 1067, 1164, 1261, 1358, 1455, 1552, 1649, 1746, 1843, 1940, 2037, 2134, 2231, 2328, 2425, 2522, 2619, 2716, 2813, 2910, 3007, 3104, 3201, 3298, 3395, 3492, 3589, 3686, 3783, 3880, 3977, 4074, 4171, 4268, 4365, 4462, 4559, 4656, 4753, 4850, 4947, 5044, 5141, 5238, 5335, 5432, 5529, 5626, 5723, 5820, 5917, 6014, 6111, 6208, 6305, 6402, 6499, 6596, 6693, 6790, 6887, 6984, 7081, 7178, 7275, 7372, 7469, 7566, 7663, 7760, 7857, 7954, 8051, 8148, 8245, 8342, 8439, 8536, 8633, 8730, 8827, 8924, 9021, 9118, 9215, 9312, 9409, 9506, 9603, 9700, 9797, 9894, 9991, 10088, 10185, 10282, 10379, 10476, 10573, 10670, 10767, 10864, 10961, 11058, 11155, 11252, 11349, 11446, 11543, 11640, 11737, 11834, 11931, 12028, 12125, 12222, 12319, 12416, 12513, 12610, 12707, 12804, 12901, 12998, 13095, 13192, 13289, 13386, 13483, 13580, 13677, 13774, 13871, 13968, 14065, 14162, 14259, 14356, 14453, 14550, 14647, 14744, 14841, 14938, 15035, 15132, 15229, 15326, 15423, 15520, 15617, 15714, 15811, 15908, 16005, 16102, 16199, 16296, 16393, 16490, 16587, 16684, 16781, 16878, 16975, 17072, 17169, 17266, 17363, 17460, 17557, 17654, 17751, 17848, 17945, 18042, 18139, 18236, 18333, 18430, 18527, 18624, 18721, 18818, 18915, 19012, 19109, 19206, 19303, 19400, 19497, 19594, 19691, 19788, 19885, 19982, 20079, 20176, 20273, 20370, 20467, 20564, 20661, 20758, 20855, 20952, 21049, 21146, 21243, 21340, 21437, 21534, 21631, 21728, 21825, 21922, 22019, 22116, 22213, 22310, 22407, 22504, 22601, 22698, 22795, 22892, 22989, 23086, 23183, 23280, 23377, 23474, 23571, 23668, 23765, 23862, 23959, 24056, 24153, 24250, 24347, 24444, 24541, 24638, 24735, 
0, 98, 196, 294, 392, 490, 588, 686, 784, 882, 980, 1078, 1176, 1274, 1372, 1470, 1568, 1666, 1764, 1862, 1960, 2058, 2156, 2254, 2352, 2450, 2548, 2646, 2744, 2842, 2940, 3038, 3136, 3234, 3332, 3430, 3528, 3626, 3724, 3822, 3920, 4018, 4116, 4214, 4312, 4410, 4508, 4606, 4704, 4802, 4900, 4998, 5096, 5194, 5292, 5390, 5488, 5586, 5684, 5782, 5880, 5978, 6076, 6174, 6272, 6370, 6468, 6566, 6664, 6762, 6860, 6958, 7056, 7154, 7252, 7350, 7448, 7546, 7644, 7742, 7840, 7938, 8036, 8134, 8232, 8330, 8428, 8526, 8624, 8722, 8820, 8918, 9016, 9114, 9212, 9310, 9408, 9506, 9604, 9702, 9800, 9898, 9996, 10094, 10192, 10290, 10388, 10486, 10584, 10682, 10780, 10878, 10976, 11074, 11172, 11270, 11368, 11466, 11564, 11662, 11760, 11858, 11956, 12054, 12152, 12250, 12348, 12446, 12544, 12642, 12740, 12838, 12936, 13034, 13132, 13230, 13328, 13426, 13524, 13622, 13720, 13818, 13916, 14014, 14112, 14210, 14308, 14406, 14504, 14602, 14700, 14798, 14896, 14994, 15092, 15190, 15288, 15386, 15484, 15582, 15680, 15778, 15876, 15974, 16072, 16170, 16268, 16366, 16464, 16562, 16660, 16758, 16856, 16954, 17052, 17150, 17248, 17346, 17444, 17542, 17640, 17738, 17836, 17934, 18032, 18130, 18228, 18326, 18424, 18522, 18620, 18718, 18816, 18914, 19012, 19110, 19208, 19306, 19404, 19502, 19600, 19698, 19796, 19894, 19992, 20090, 20188, 20286, 20384, 20482, 20580, 20678, 20776, 20874, 20972, 21070, 21168, 21266, 21364, 21462, 21560, 21658, 21756, 21854, 21952, 22050, 22148, 22246, 22344, 22442, 22540, 22638, 22736, 22834, 22932, 23030, 23128, 23226, 23324, 23422, 23520, 23618, 23716, 23814, 23912, 24010, 24108, 24206, 24304, 24402, 24500, 24598, 24696, 24794, 24892, 24990, 
0, 99, 198, 297, 396, 495, 594, 693, 792, 891, 990, 1089, 1188, 1287, 1386, 1485, 1584, 1683, 1782, 1881, 1980, 2079, 2178, 2277, 2376, 2475, 2574, 2673, 2772, 2871, 2970, 3069, 3168, 3267, 3366, 3465, 3564, 3663, 3762, 3861, 3960, 4059, 4158, 4257, 4356, 4455, 4554, 4653, 4752, 4851, 4950, 5049, 5148, 5247, 5346, 5445, 5544, 5643, 5742, 5841, 5940, 6039, 6138, 6237, 6336, 6435, 6534, 6633, 6732, 6831, 6930, 7029, 7128, 7227, 7326, 7425, 7524, 7623, 7722, 7821, 7920, 8019, 8118, 8217, 8316, 8415, 8514, 8613, 8712, 8811, 8910, 9009, 9108, 9207, 9306, 9405, 9504, 9603, 9702, 9801, 9900, 9999, 10098, 10197, 10296, 10395, 10494, 10593, 10692, 10791, 10890, 10989, 11088, 11187, 11286, 11385, 11484, 11583, 11682, 11781, 11880, 11979, 12078, 12177, 12276, 12375, 12474, 12573, 12672, 12771, 12870, 12969, 13068, 13167, 13266, 13365, 13464, 13563, 13662, 13761, 13860, 13959, 14058, 14157, 14256, 14355, 14454, 14553, 14652, 14751, 14850, 14949, 15048, 15147, 15246, 15345, 15444, 15543, 15642, 15741, 15840, 15939, 16038, 16137, 16236, 16335, 16434, 16533, 16632, 16731, 16830, 16929, 17028, 17127, 17226, 17325, 17424, 17523, 17622, 17721, 17820, 17919, 18018, 18117, 18216, 18315, 18414, 18513, 18612, 18711, 18810, 18909, 19008, 19107, 19206, 19305, 19404, 19503, 19602, 19701, 19800, 19899, 19998, 20097, 20196, 20295, 20394, 20493, 20592, 20691, 20790, 20889, 20988, 21087, 21186, 21285, 21384, 21483, 21582, 21681, 21780, 21879, 21978, 22077, 22176, 22275, 22374, 22473, 22572, 22671, 22770, 22869, 22968, 23067, 23166, 23265, 23364, 23463, 23562, 23661, 23760, 23859, 23958, 24057, 24156, 24255, 24354, 24453, 24552, 24651, 24750, 24849, 24948, 25047, 25146, 25245, 
0, 100, 200, 300, 400, 500, 600, 700, 800, 900, 1000, 1100, 1200, 1300, 1400, 1500, 1600, 1700, 1800, 1900, 2000, 2100, 2200, 2300, 2400, 2500, 2600, 2700, 2800, 2900, 3000, 3100, 3200, 3300, 3400, 3500, 3600, 3700, 3800, 3900, 4000, 4100, 4200, 4300, 4400, 4500, 4600, 4700, 4800, 4900, 5000, 5100, 5200, 5300, 5400, 5500, 5600, 5700, 5800, 5900, 6000, 6100, 6200, 6300, 6400, 6500, 6600, 6700, 6800, 6900, 7000, 7100, 7200, 7300, 7400, 7500, 7600, 7700, 7800, 7900, 8000, 8100, 8200, 8300, 8400, 8500, 8600, 8700, 8800, 8900, 9000, 9100, 9200, 9300, 9400, 9500, 9600, 9700, 9800, 9900, 10000, 10100, 10200, 10300, 10400, 10500, 10600, 10700, 10800, 10900, 11000, 11100, 11200, 11300, 11400, 11500, 11600, 11700, 11800, 11900, 12000, 12100, 12200, 12300, 12400, 12500, 12600, 12700, 12800, 12900, 13000, 13100, 13200, 13300, 13400, 13500, 13600, 13700, 13800, 13900, 14000, 14100, 14200, 14300, 14400, 14500, 14600, 14700, 14800, 14900, 15000, 15100, 15200, 15300, 15400, 15500, 15600, 15700, 15800, 15900, 16000, 16100, 16200, 16300, 16400, 16500, 16600, 16700, 16800, 16900, 17000, 17100, 17200, 17300, 17400, 17500, 17600, 17700, 17800, 17900, 18000, 18100, 18200, 18300, 18400, 18500, 18600, 18700, 18800, 18900, 19000, 19100, 19200, 19300, 19400, 19500, 19600, 19700, 19800, 19900, 20000, 20100, 20200, 20300, 20400, 20500, 20600, 20700, 20800, 20900, 21000, 21100, 21200, 21300, 21400, 21500, 21600, 21700, 21800, 21900, 22000, 22100, 22200, 22300, 22400, 22500, 22600, 22700, 22800, 22900, 23000, 23100, 23200, 23300, 23400, 23500, 23600, 23700, 23800, 23900, 24000, 24100, 24200, 24300, 24400, 24500, 24600, 24700, 24800, 24900, 25000, 25100, 25200, 25300, 25400, 25500, 
0, 101, 202, 303, 404, 505, 606, 707, 808, 909, 1010, 1111, 1212, 1313, 1414, 1515, 1616, 1717, 1818, 1919, 2020, 2121, 2222, 2323, 2424, 2525, 2626, 2727, 2828, 2929, 3030, 3131, 3232, 3333, 3434, 3535, 3636, 3737, 3838, 3939, 4040, 4141, 4242, 4343, 4444, 4545, 4646, 4747, 4848, 4949, 5050, 5151, 5252, 5353, 5454, 5555, 5656, 5757, 5858, 5959, 6060, 6161, 6262, 6363, 6464, 6565, 6666, 6767, 6868, 6969, 7070, 7171, 7272, 7373, 7474, 7575, 7676, 7777, 7878, 7979, 8080, 8181, 8282, 8383, 8484, 8585, 8686, 8787, 8888, 8989, 9090, 9191, 9292, 9393, 9494, 9595, 9696, 9797, 9898, 9999, 10100, 10201, 10302, 10403, 10504, 10605, 10706, 10807, 10908, 11009, 11110, 11211, 11312, 11413, 11514, 11615, 11716, 11817, 11918, 12019, 12120, 12221, 12322, 12423, 12524, 12625, 12726, 12827, 12928, 13029, 13130, 13231, 13332, 13433, 13534, 13635, 13736, 13837, 13938, 14039, 14140, 14241, 14342, 14443, 14544, 14645, 14746, 14847, 14948, 15049, 15150, 15251, 15352, 15453, 15554, 15655, 15756, 15857, 15958, 16059, 16160, 16261, 16362, 16463, 16564, 16665, 16766, 16867, 16968, 17069, 17170, 17271, 17372, 17473, 17574, 17675, 17776, 17877, 17978, 18079, 18180, 18281, 18382, 18483, 18584, 18685, 18786, 18887, 18988, 19089, 19190, 19291, 19392, 19493, 19594, 19695, 19796, 19897, 19998, 20099, 20200, 20301, 20402, 20503, 20604, 20705, 20806, 20907, 21008, 21109, 21210, 21311, 21412, 21513, 21614, 21715, 21816, 21917, 22018, 22119, 22220, 22321, 22422, 22523, 22624, 22725, 22826, 22927, 23028, 23129, 23230, 23331, 23432, 23533, 23634, 23735, 23836, 23937, 24038, 24139, 24240, 24341, 24442, 24543, 24644, 24745, 24846, 24947, 25048, 25149, 25250, 25351, 25452, 25553, 25654, 25755, 
0, 102, 204, 306, 408, 510, 612, 714, 816, 918, 1020, 1122, 1224, 1326, 1428, 1530, 1632, 1734, 1836, 1938, 2040, 2142, 2244, 2346, 2448, 2550, 2652, 2754, 2856, 2958, 3060, 3162, 3264, 3366, 3468, 3570, 3672, 3774, 3876, 3978, 4080, 4182, 4284, 4386, 4488, 4590, 4692, 4794, 4896, 4998, 5100, 5202, 5304, 5406, 5508, 5610, 5712, 5814, 5916, 6018, 6120, 6222, 6324, 6426, 6528, 6630, 6732, 6834, 6936, 7038, 7140, 7242, 7344, 7446, 7548, 7650, 7752, 7854, 7956, 8058, 8160, 8262, 8364, 8466, 8568, 8670, 8772, 8874, 8976, 9078, 9180, 9282, 9384, 9486, 9588, 9690, 9792, 9894, 9996, 10098, 10200, 10302, 10404, 10506, 10608, 10710, 10812, 10914, 11016, 11118, 11220, 11322, 11424, 11526, 11628, 11730, 11832, 11934, 12036, 12138, 12240, 12342, 12444, 12546, 12648, 12750, 12852, 12954, 13056, 13158, 13260, 13362, 13464, 13566, 13668, 13770, 13872, 13974, 14076, 14178, 14280, 14382, 14484, 14586, 14688, 14790, 14892, 14994, 15096, 15198, 15300, 15402, 15504, 15606, 15708, 15810, 15912, 16014, 16116, 16218, 16320, 16422, 16524, 16626, 16728, 16830, 16932, 17034, 17136, 17238, 17340, 17442, 17544, 17646, 17748, 17850, 17952, 18054, 18156, 18258, 18360, 18462, 18564, 18666, 18768, 18870, 18972, 19074, 19176, 19278, 19380, 19482, 19584, 19686, 19788, 19890, 19992, 20094, 20196, 20298, 20400, 20502, 20604, 20706, 20808, 20910, 21012, 21114, 21216, 21318, 21420, 21522, 21624, 21726, 21828, 21930, 22032, 22134, 22236, 22338, 22440, 22542, 22644, 22746, 22848, 22950, 23052, 23154, 23256, 23358, 23460, 23562, 23664, 23766, 23868, 23970, 24072, 24174, 24276, 24378, 24480, 24582, 24684, 24786, 24888, 24990, 25092, 25194, 25296, 25398, 25500, 25602, 25704, 25806, 25908, 26010, 
0, 103, 206, 309, 412, 515, 618, 721, 824, 927, 1030, 1133, 1236, 1339, 1442, 1545, 1648, 1751, 1854, 1957, 2060, 2163, 2266, 2369, 2472, 2575, 2678, 2781, 2884, 2987, 3090, 3193, 3296, 3399, 3502, 3605, 3708, 3811, 3914, 4017, 4120, 4223, 4326, 4429, 4532, 4635, 4738, 4841, 4944, 5047, 5150, 5253, 5356, 5459, 5562, 5665, 5768, 5871, 5974, 6077, 6180, 6283, 6386, 6489, 6592, 6695, 6798, 6901, 7004, 7107, 7210, 7313, 7416, 7519, 7622, 7725, 7828, 7931, 8034, 8137, 8240, 8343, 8446, 8549, 8652, 8755, 8858, 8961, 9064, 9167, 9270, 9373, 9476, 9579, 9682, 9785, 9888, 9991, 10094, 10197, 10300, 10403, 10506, 10609, 10712, 10815, 10918, 11021, 11124, 11227, 11330, 11433, 11536, 11639, 11742, 11845, 11948, 12051, 12154, 12257, 12360, 12463, 12566, 12669, 12772, 12875, 12978, 13081, 13184, 13287, 13390, 13493, 13596, 13699, 13802, 13905, 14008, 14111, 14214, 14317, 14420, 14523, 14626, 14729, 14832, 14935, 15038, 15141, 15244, 15347, 15450, 15553, 15656, 15759, 15862, 15965, 16068, 16171, 16274, 16377, 16480, 16583, 16686, 16789, 16892, 16995, 17098, 17201, 17304, 17407, 17510, 17613, 17716, 17819, 17922, 18025, 18128, 18231, 18334, 18437, 18540, 18643, 18746, 18849, 18952, 19055, 19158, 19261, 19364, 19467, 19570, 19673, 19776, 19879, 19982, 20085, 20188, 20291, 20394, 20497, 20600, 20703, 20806, 20909, 21012, 21115, 21218, 21321, 21424, 21527, 21630, 21733, 21836, 21939, 22042, 22145, 22248, 22351, 22454, 22557, 22660, 22763, 22866, 22969, 23072, 23175, 23278, 23381, 23484, 23587, 23690, 23793, 23896, 23999, 24102, 24205, 24308, 24411, 24514, 24617, 24720, 24823, 24926, 25029, 25132, 25235, 25338, 25441, 25544, 25647, 25750, 25853, 25956, 26059, 26162, 26265, 
0, 104, 208, 312, 416, 520, 624, 728, 832, 936, 1040, 1144, 1248, 1352, 1456, 1560, 1664, 1768, 1872, 1976, 2080, 2184, 2288, 2392, 2496, 2600, 2704, 2808, 2912, 3016, 3120, 3224, 3328, 3432, 3536, 3640, 3744, 3848, 3952, 4056, 4160, 4264, 4368, 4472, 4576, 4680, 4784, 4888, 4992, 5096, 5200, 5304, 5408, 5512, 5616, 5720, 5824, 5928, 6032, 6136, 6240, 6344, 6448, 6552, 6656, 6760, 6864, 6968, 7072, 7176, 7280, 7384, 7488, 7592, 7696, 7800, 7904, 8008, 8112, 8216, 8320, 8424, 8528, 8632, 8736, 8840, 8944, 9048, 9152, 9256, 9360, 9464, 9568, 9672, 9776, 9880, 9984, 10088, 10192, 10296, 10400, 10504, 10608, 10712, 10816, 10920, 11024, 11128, 11232, 11336, 11440, 11544, 11648, 11752, 11856, 11960, 12064, 12168, 12272, 12376, 12480, 12584, 12688, 12792, 12896, 13000, 13104, 13208, 13312, 13416, 13520, 13624, 13728, 13832, 13936, 14040, 14144, 14248, 14352, 14456, 14560, 14664, 14768, 14872, 14976, 15080, 15184, 15288, 15392, 15496, 15600, 15704, 15808, 15912, 16016, 16120, 16224, 16328, 16432, 16536, 16640, 16744, 16848, 16952, 17056, 17160, 17264, 17368, 17472, 17576, 17680, 17784, 17888, 17992, 18096, 18200, 18304, 18408, 18512, 18616, 18720, 18824, 18928, 19032, 19136, 19240, 19344, 19448, 19552, 19656, 19760, 19864, 19968, 20072, 20176, 20280, 20384, 20488, 20592, 20696, 20800, 20904, 21008, 21112, 21216, 21320, 21424, 21528, 21632, 21736, 21840, 21944, 22048, 22152, 22256, 22360, 22464, 22568, 22672, 22776, 22880, 22984, 23088, 23192, 23296, 23400, 23504, 23608, 23712, 23816, 23920, 24024, 24128, 24232, 24336, 24440, 24544, 24648, 24752, 24856, 24960, 25064, 25168, 25272, 25376, 25480, 25584, 25688, 25792, 25896, 26000, 26104, 26208, 26312, 26416, 26520, 
0, 105, 210, 315, 420, 525, 630, 735, 840, 945, 1050, 1155, 1260, 1365, 1470, 1575, 1680, 1785, 1890, 1995, 2100, 2205, 2310, 2415, 2520, 2625, 2730, 2835, 2940, 3045, 3150, 3255, 3360, 3465, 3570, 3675, 3780, 3885, 3990, 4095, 4200, 4305, 4410, 4515, 4620, 4725, 4830, 4935, 5040, 5145, 5250, 5355, 5460, 5565, 5670, 5775, 5880, 5985, 6090, 6195, 6300, 6405, 6510, 6615, 6720, 6825, 6930, 7035, 7140, 7245, 7350, 7455, 7560, 7665, 7770, 7875, 7980, 8085, 8190, 8295, 8400, 8505, 8610, 8715, 8820, 8925, 9030, 9135, 9240, 9345, 9450, 9555, 9660, 9765, 9870, 9975, 10080, 10185, 10290, 10395, 10500, 10605, 10710, 10815, 10920, 11025, 11130, 11235, 11340, 11445, 11550, 11655, 11760, 11865, 11970, 12075, 12180, 12285, 12390, 12495, 12600, 12705, 12810, 12915, 13020, 13125, 13230, 13335, 13440, 13545, 13650, 13755, 13860, 13965, 14070, 14175, 14280, 14385, 14490, 14595, 14700, 14805, 14910, 15015, 15120, 15225, 15330, 15435, 15540, 15645, 15750, 15855, 15960, 16065, 16170, 16275, 16380, 16485, 16590, 16695, 16800, 16905, 17010, 17115, 17220, 17325, 17430, 17535, 17640, 17745, 17850, 17955, 18060, 18165, 18270, 18375, 18480, 18585, 18690, 18795, 18900, 19005, 19110, 19215, 19320, 19425, 19530, 19635, 19740, 19845, 19950, 20055, 20160, 20265, 20370, 20475, 20580, 20685, 20790, 20895, 21000, 21105, 21210, 21315, 21420, 21525, 21630, 21735, 21840, 21945, 22050, 22155, 22260, 22365, 22470, 22575, 22680, 22785, 22890, 22995, 23100, 23205, 23310, 23415, 23520, 23625, 23730, 23835, 23940, 24045, 24150, 24255, 24360, 24465, 24570, 24675, 24780, 24885, 24990, 25095, 25200, 25305, 25410, 25515, 25620, 25725, 25830, 25935, 26040, 26145, 26250, 26355, 26460, 26565, 26670, 26775, 
0, 106, 212, 318, 424, 530, 636, 742, 848, 954, 1060, 1166, 1272, 1378, 1484, 1590, 1696, 1802, 1908, 2014, 2120, 2226, 2332, 2438, 2544, 2650, 2756, 2862, 2968, 3074, 3180, 3286, 3392, 3498, 3604, 3710, 3816, 3922, 4028, 4134, 4240, 4346, 4452, 4558, 4664, 4770, 4876, 4982, 5088, 5194, 5300, 5406, 5512, 5618, 5724, 5830, 5936, 6042, 6148, 6254, 6360, 6466, 6572, 6678, 6784, 6890, 6996, 7102, 7208, 7314, 7420, 7526, 7632, 7738, 7844, 7950, 8056, 8162, 8268, 8374, 8480, 8586, 8692, 8798, 8904, 9010, 9116, 9222, 9328, 9434, 9540, 9646, 9752, 9858, 9964, 10070, 10176, 10282, 10388, 10494, 10600, 10706, 10812, 10918, 11024, 11130, 11236, 11342, 11448, 11554, 11660, 11766, 11872, 11978, 12084, 12190, 12296, 12402, 12508, 12614, 12720, 12826, 12932, 13038, 13144, 13250, 13356, 13462, 13568, 13674, 13780, 13886, 13992, 14098, 14204, 14310, 14416, 14522, 14628, 14734, 14840, 14946, 15052, 15158, 15264, 15370, 15476, 15582, 15688, 15794, 15900, 16006, 16112, 16218, 16324, 16430, 16536, 16642, 16748, 16854, 16960, 17066, 17172, 17278, 17384, 17490, 17596, 17702, 17808, 17914, 18020, 18126, 18232, 18338, 18444, 18550, 18656, 18762, 18868, 18974, 19080, 19186, 19292, 19398, 19504, 19610, 19716, 19822, 19928, 20034, 20140, 20246, 20352, 20458, 20564, 20670, 20776, 20882, 20988, 21094, 21200, 21306, 21412, 21518, 21624, 21730, 21836, 21942, 22048, 22154, 22260, 22366, 22472, 22578, 22684, 22790, 22896, 23002, 23108, 23214, 23320, 23426, 23532, 23638, 23744, 23850, 23956, 24062, 24168, 24274, 24380, 24486, 24592, 24698, 24804, 24910, 25016, 25122, 25228, 25334, 25440, 25546, 25652, 25758, 25864, 25970, 26076, 26182, 26288, 26394, 26500, 26606, 26712, 26818, 26924, 27030, 
0, 107, 214, 321, 428, 535, 642, 749, 856, 963, 1070, 1177, 1284, 1391, 1498, 1605, 1712, 1819, 1926, 2033, 2140, 2247, 2354, 2461, 2568, 2675, 2782, 2889, 2996, 3103, 3210, 3317, 3424, 3531, 3638, 3745, 3852, 3959, 4066, 4173, 4280, 4387, 4494, 4601, 4708, 4815, 4922, 5029, 5136, 5243, 5350, 5457, 5564, 5671, 5778, 5885, 5992, 6099, 6206, 6313, 6420, 6527, 6634, 6741, 6848, 6955, 7062, 7169, 7276, 7383, 7490, 7597, 7704, 7811, 7918, 8025, 8132, 8239, 8346, 8453, 8560, 8667, 8774, 8881, 8988, 9095, 9202, 9309, 9416, 9523, 9630, 9737, 9844, 9951, 10058, 10165, 10272, 10379, 10486, 10593, 10700, 10807, 10914, 11021, 11128, 11235, 11342, 11449, 11556, 11663, 11770, 11877, 11984, 12091, 12198, 12305, 12412, 12519, 12626, 12733, 12840, 12947, 13054, 13161, 13268, 13375, 13482, 13589, 13696, 13803, 13910, 14017, 14124, 14231, 14338, 14445, 14552, 14659, 14766, 14873, 14980, 15087, 15194, 15301, 15408, 15515, 15622, 15729, 15836, 15943, 16050, 16157, 16264, 16371, 16478, 16585, 16692, 16799, 16906, 17013, 17120, 17227, 17334, 17441, 17548, 17655, 17762, 17869, 17976, 18083, 18190, 18297, 18404, 18511, 18618, 18725, 18832, 18939, 19046, 19153, 19260, 19367, 19474, 19581, 19688, 19795, 19902, 20009, 20116, 20223, 20330, 20437, 20544, 20651, 20758, 20865, 20972, 21079, 21186, 21293, 21400, 21507, 21614, 21721, 21828, 21935, 22042, 22149, 22256, 22363, 22470, 22577, 22684, 22791, 22898, 23005, 23112, 23219, 23326, 23433, 23540, 23647, 23754, 23861, 23968, 24075, 24182, 24289, 24396, 24503, 24610, 24717, 24824, 24931, 25038, 25145, 25252, 25359, 25466, 25573, 25680, 25787, 25894, 26001, 26108, 26215, 26322, 26429, 26536, 26643, 26750, 26857, 26964, 27071, 27178, 27285, 
0, 108, 216, 324, 432, 540, 648, 756, 864, 972, 1080, 1188, 1296, 1404, 1512, 1620, 1728, 1836, 1944, 2052, 2160, 2268, 2376, 2484, 2592, 2700, 2808, 2916, 3024, 3132, 3240, 3348, 3456, 3564, 3672, 3780, 3888, 3996, 4104, 4212, 4320, 4428, 4536, 4644, 4752, 4860, 4968, 5076, 5184, 5292, 5400, 5508, 5616, 5724, 5832, 5940, 6048, 6156, 6264, 6372, 6480, 6588, 6696, 6804, 6912, 7020, 7128, 7236, 7344, 7452, 7560, 7668, 7776, 7884, 7992, 8100, 8208, 8316, 8424, 8532, 8640, 8748, 8856, 8964, 9072, 9180, 9288, 9396, 9504, 9612, 9720, 9828, 9936, 10044, 10152, 10260, 10368, 10476, 10584, 10692, 10800, 10908, 11016, 11124, 11232, 11340, 11448, 11556, 11664, 11772, 11880, 11988, 12096, 12204, 12312, 12420, 12528, 12636, 12744, 12852, 12960, 13068, 13176, 13284, 13392, 13500, 13608, 13716, 13824, 13932, 14040, 14148, 14256, 14364, 14472, 14580, 14688, 14796, 14904, 15012, 15120, 15228, 15336, 15444, 15552, 15660, 15768, 15876, 15984, 16092, 16200, 16308, 16416, 16524, 16632, 16740, 16848, 16956, 17064, 17172, 17280, 17388, 17496, 17604, 17712, 17820, 17928, 18036, 18144, 18252, 18360, 18468, 18576, 18684, 18792, 18900, 19008, 19116, 19224, 19332, 19440, 19548, 19656, 19764, 19872, 19980, 20088, 20196, 20304, 20412, 20520, 20628, 20736, 20844, 20952, 21060, 21168, 21276, 21384, 21492, 21600, 21708, 21816, 21924, 22032, 22140, 22248, 22356, 22464, 22572, 22680, 22788, 22896, 23004, 23112, 23220, 23328, 23436, 23544, 23652, 23760, 23868, 23976, 24084, 24192, 24300, 24408, 24516, 24624, 24732, 24840, 24948, 25056, 25164, 25272, 25380, 25488, 25596, 25704, 25812, 25920, 26028, 26136, 26244, 26352, 26460, 26568, 26676, 26784, 26892, 27000, 27108, 27216, 27324, 27432, 27540, 
0, 109, 218, 327, 436, 545, 654, 763, 872, 981, 1090, 1199, 1308, 1417, 1526, 1635, 1744, 1853, 1962, 2071, 2180, 2289, 2398, 2507, 2616, 2725, 2834, 2943, 3052, 3161, 3270, 3379, 3488, 3597, 3706, 3815, 3924, 4033, 4142, 4251, 4360, 4469, 4578, 4687, 4796, 4905, 5014, 5123, 5232, 5341, 5450, 5559, 5668, 5777, 5886, 5995, 6104, 6213, 6322, 6431, 6540, 6649, 6758, 6867, 6976, 7085, 7194, 7303, 7412, 7521, 7630, 7739, 7848, 7957, 8066, 8175, 8284, 8393, 8502, 8611, 8720, 8829, 8938, 9047, 9156, 9265, 9374, 9483, 9592, 9701, 9810, 9919, 10028, 10137, 10246, 10355, 10464, 10573, 10682, 10791, 10900, 11009, 11118, 11227, 11336, 11445, 11554, 11663, 11772, 11881, 11990, 12099, 12208, 12317, 12426, 12535, 12644, 12753, 12862, 12971, 13080, 13189, 13298, 13407, 13516, 13625, 13734, 13843, 13952, 14061, 14170, 14279, 14388, 14497, 14606, 14715, 14824, 14933, 15042, 15151, 15260, 15369, 15478, 15587, 15696, 15805, 15914, 16023, 16132, 16241, 16350, 16459, 16568, 16677, 16786, 16895, 17004, 17113, 17222, 17331, 17440, 17549, 17658, 17767, 17876, 17985, 18094, 18203, 18312, 18421, 18530, 18639, 18748, 18857, 18966, 19075, 19184, 19293, 19402, 19511, 19620, 19729, 19838, 19947, 20056, 20165, 20274, 20383, 20492, 20601, 20710, 20819, 20928, 21037, 21146, 21255, 21364, 21473, 21582, 21691, 21800, 21909, 22018, 22127, 22236, 22345, 22454, 22563, 22672, 22781, 22890, 22999, 23108, 23217, 23326, 23435, 23544, 23653, 23762, 23871, 23980, 24089, 24198, 24307, 24416, 24525, 24634, 24743, 24852, 24961, 25070, 25179, 25288, 25397, 25506, 25615, 25724, 25833, 25942, 26051, 26160, 26269, 26378, 26487, 26596, 26705, 26814, 26923, 27032, 27141, 27250, 27359, 27468, 27577, 27686, 27795, 
0, 110, 220, 330, 440, 550, 660, 770, 880, 990, 1100, 1210, 1320, 1430, 1540, 1650, 1760, 1870, 1980, 2090, 2200, 2310, 2420, 2530, 2640, 2750, 2860, 2970, 3080, 3190, 3300, 3410, 3520, 3630, 3740, 3850, 3960, 4070, 4180, 4290, 4400, 4510, 4620, 4730, 4840, 4950, 5060, 5170, 5280, 5390, 5500, 5610, 5720, 5830, 5940, 6050, 6160, 6270, 6380, 6490, 6600, 6710, 6820, 6930, 7040, 7150, 7260, 7370, 7480, 7590, 7700, 7810, 7920, 8030, 8140, 8250, 8360, 8470, 8580, 8690, 8800, 8910, 9020, 9130, 9240, 9350, 9460, 9570, 9680, 9790, 9900, 10010, 10120, 10230, 10340, 10450, 10560, 10670, 10780, 10890, 11000, 11110, 11220, 11330, 11440, 11550, 11660, 11770, 11880, 11990, 12100, 12210, 12320, 12430, 12540, 12650, 12760, 12870, 12980, 13090, 13200, 13310, 13420, 13530, 13640, 13750, 13860, 13970, 14080, 14190, 14300, 14410, 14520, 14630, 14740, 14850, 14960, 15070, 15180, 15290, 15400, 15510, 15620, 15730, 15840, 15950, 16060, 16170, 16280, 16390, 16500, 16610, 16720, 16830, 16940, 17050, 17160, 17270, 17380, 17490, 17600, 17710, 17820, 17930, 18040, 18150, 18260, 18370, 18480, 18590, 18700, 18810, 18920, 19030, 19140, 19250, 19360, 19470, 19580, 19690, 19800, 19910, 20020, 20130, 20240, 20350, 20460, 20570, 20680, 20790, 20900, 21010, 21120, 21230, 21340, 21450, 21560, 21670, 21780, 21890, 22000, 22110, 22220, 22330, 22440, 22550, 22660, 22770, 22880, 22990, 23100, 23210, 23320, 23430, 23540, 23650, 23760, 23870, 23980, 24090, 24200, 24310, 24420, 24530, 24640, 24750, 24860, 24970, 25080, 25190, 25300, 25410, 25520, 25630, 25740, 25850, 25960, 26070, 26180, 26290, 26400, 26510, 26620, 26730, 26840, 26950, 27060, 27170, 27280, 27390, 27500, 27610, 27720, 27830, 27940, 28050, 
0, 111, 222, 333, 444, 555, 666, 777, 888, 999, 1110, 1221, 1332, 1443, 1554, 1665, 1776, 1887, 1998, 2109, 2220, 2331, 2442, 2553, 2664, 2775, 2886, 2997, 3108, 3219, 3330, 3441, 3552, 3663, 3774, 3885, 3996, 4107, 4218, 4329, 4440, 4551, 4662, 4773, 4884, 4995, 5106, 5217, 5328, 5439, 5550, 5661, 5772, 5883, 5994, 6105, 6216, 6327, 6438, 6549, 6660, 6771, 6882, 6993, 7104, 7215, 7326, 7437, 7548, 7659, 7770, 7881, 7992, 8103, 8214, 8325, 8436, 8547, 8658, 8769, 8880, 8991, 9102, 9213, 9324, 9435, 9546, 9657, 9768, 9879, 9990, 10101, 10212, 10323, 10434, 10545, 10656, 10767, 10878, 10989, 11100, 11211, 11322, 11433, 11544, 11655, 11766, 11877, 11988, 12099, 12210, 12321, 12432, 12543, 12654, 12765, 12876, 12987, 13098, 13209, 13320, 13431, 13542, 13653, 13764, 13875, 13986, 14097, 14208, 14319, 14430, 14541, 14652, 14763, 14874, 14985, 15096, 15207, 15318, 15429, 15540, 15651, 15762, 15873, 15984, 16095, 16206, 16317, 16428, 16539, 16650, 16761, 16872, 16983, 17094, 17205, 17316, 17427, 17538, 17649, 17760, 17871, 17982, 18093, 18204, 18315, 18426, 18537, 18648, 18759, 18870, 18981, 19092, 19203, 19314, 19425, 19536, 19647, 19758, 19869, 19980, 20091, 20202, 20313, 20424, 20535, 20646, 20757, 20868, 20979, 21090, 21201, 21312, 21423, 21534, 21645, 21756, 21867, 21978, 22089, 22200, 22311, 22422, 22533, 22644, 22755, 22866, 22977, 23088, 23199, 23310, 23421, 23532, 23643, 23754, 23865, 23976, 24087, 24198, 24309, 24420, 24531, 24642, 24753, 24864, 24975, 25086, 25197, 25308, 25419, 25530, 25641, 25752, 25863, 25974, 26085, 26196, 26307, 26418, 26529, 26640, 26751, 26862, 26973, 27084, 27195, 27306, 27417, 27528, 27639, 27750, 27861, 27972, 28083, 28194, 28305, 
0, 112, 224, 336, 448, 560, 672, 784, 896, 1008, 1120, 1232, 1344, 1456, 1568, 1680, 1792, 1904, 2016, 2128, 2240, 2352, 2464, 2576, 2688, 2800, 2912, 3024, 3136, 3248, 3360, 3472, 3584, 3696, 3808, 3920, 4032, 4144, 4256, 4368, 4480, 4592, 4704, 4816, 4928, 5040, 5152, 5264, 5376, 5488, 5600, 5712, 5824, 5936, 6048, 6160, 6272, 6384, 6496, 6608, 6720, 6832, 6944, 7056, 7168, 7280, 7392, 7504, 7616, 7728, 7840, 7952, 8064, 8176, 8288, 8400, 8512, 8624, 8736, 8848, 8960, 9072, 9184, 9296, 9408, 9520, 9632, 9744, 9856, 9968, 10080, 10192, 10304, 10416, 10528, 10640, 10752, 10864, 10976, 11088, 11200, 11312, 11424, 11536, 11648, 11760, 11872, 11984, 12096, 12208, 12320, 12432, 12544, 12656, 12768, 12880, 12992, 13104, 13216, 13328, 13440, 13552, 13664, 13776, 13888, 14000, 14112, 14224, 14336, 14448, 14560, 14672, 14784, 14896, 15008, 15120, 15232, 15344, 15456, 15568, 15680, 15792, 15904, 16016, 16128, 16240, 16352, 16464, 16576, 16688, 16800, 16912, 17024, 17136, 17248, 17360, 17472, 17584, 17696, 17808, 17920, 18032, 18144, 18256, 18368, 18480, 18592, 18704, 18816, 18928, 19040, 19152, 19264, 19376, 19488, 19600, 19712, 19824, 19936, 20048, 20160, 20272, 20384, 20496, 20608, 20720, 20832, 20944, 21056, 21168, 21280, 21392, 21504, 21616, 21728, 21840, 21952, 22064, 22176, 22288, 22400, 22512, 22624, 22736, 22848, 22960, 23072, 23184, 23296, 23408, 23520, 23632, 23744, 23856, 23968, 24080, 24192, 24304, 24416, 24528, 24640, 24752, 24864, 24976, 25088, 25200, 25312, 25424, 25536, 25648, 25760, 25872, 25984, 26096, 26208, 26320, 26432, 26544, 26656, 26768, 26880, 26992, 27104, 27216, 27328, 27440, 27552, 27664, 27776, 27888, 28000, 28112, 28224, 28336, 28448, 28560, 
0, 113, 226, 339, 452, 565, 678, 791, 904, 1017, 1130, 1243, 1356, 1469, 1582, 1695, 1808, 1921, 2034, 2147, 2260, 2373, 2486, 2599, 2712, 2825, 2938, 3051, 3164, 3277, 3390, 3503, 3616, 3729, 3842, 3955, 4068, 4181, 4294, 4407, 4520, 4633, 4746, 4859, 4972, 5085, 5198, 5311, 5424, 5537, 5650, 5763, 5876, 5989, 6102, 6215, 6328, 6441, 6554, 6667, 6780, 6893, 7006, 7119, 7232, 7345, 7458, 7571, 7684, 7797, 7910, 8023, 8136, 8249, 8362, 8475, 8588, 8701, 8814, 8927, 9040, 9153, 9266, 9379, 9492, 9605, 9718, 9831, 9944, 10057, 10170, 10283, 10396, 10509, 10622, 10735, 10848, 10961, 11074, 11187, 11300, 11413, 11526, 11639, 11752, 11865, 11978, 12091, 12204, 12317, 12430, 12543, 12656, 12769, 12882, 12995, 13108, 13221, 13334, 13447, 13560, 13673, 13786, 13899, 14012, 14125, 14238, 14351, 14464, 14577, 14690, 14803, 14916, 15029, 15142, 15255, 15368, 15481, 15594, 15707, 15820, 15933, 16046, 16159, 16272, 16385, 16498, 16611, 16724, 16837, 16950, 17063, 17176, 17289, 17402, 17515, 17628, 17741, 17854, 17967, 18080, 18193, 18306, 18419, 18532, 18645, 18758, 18871, 18984, 19097, 19210, 19323, 19436, 19549, 19662, 19775, 19888, 20001, 20114, 20227, 20340, 20453, 20566, 20679, 20792, 20905, 21018, 21131, 21244, 21357, 21470, 21583, 21696, 21809, 21922, 22035, 22148, 22261, 22374, 22487, 22600, 22713, 22826, 22939, 23052, 23165, 23278, 23391, 23504, 23617, 23730, 23843, 23956, 24069, 24182, 24295, 24408, 24521, 24634, 24747, 24860, 24973, 25086, 25199, 25312, 25425, 25538, 25651, 25764, 25877, 25990, 26103, 26216, 26329, 26442, 26555, 26668, 26781, 26894, 27007, 27120, 27233, 27346, 27459, 27572, 27685, 27798, 27911, 28024, 28137, 28250, 28363, 28476, 28589, 28702, 28815, 
0, 114, 228, 342, 456, 570, 684, 798, 912, 1026, 1140, 1254, 1368, 1482, 1596, 1710, 1824, 1938, 2052, 2166, 2280, 2394, 2508, 2622, 2736, 2850, 2964, 3078, 3192, 3306, 3420, 3534, 3648, 3762, 3876, 3990, 4104, 4218, 4332, 4446, 4560, 4674, 4788, 4902, 5016, 5130, 5244, 5358, 5472, 5586, 5700, 5814, 5928, 6042, 6156, 6270, 6384, 6498, 6612, 6726, 6840, 6954, 7068, 7182, 7296, 7410, 7524, 7638, 7752, 7866, 7980, 8094, 8208, 8322, 8436, 8550, 8664, 8778, 8892, 9006, 9120, 9234, 9348, 9462, 9576, 9690, 9804, 9918, 10032, 10146, 10260, 10374, 10488, 10602, 10716, 10830, 10944, 11058, 11172, 11286, 11400, 11514, 11628, 11742, 11856, 11970, 12084, 12198, 12312, 12426, 12540, 12654, 12768, 12882, 12996, 13110, 13224, 13338, 13452, 13566, 13680, 13794, 13908, 14022, 14136, 14250, 14364, 14478, 14592, 14706, 14820, 14934, 15048, 15162, 15276, 15390, 15504, 15618, 15732, 15846, 15960, 16074, 16188, 16302, 16416, 16530, 16644, 16758, 16872, 16986, 17100, 17214, 17328, 17442, 17556, 17670, 17784, 17898, 18012, 18126, 18240, 18354, 18468, 18582, 18696, 18810, 18924, 19038, 19152, 19266, 19380, 19494, 19608, 19722, 19836, 19950, 20064, 20178, 20292, 20406, 20520, 20634, 20748, 20862, 20976, 21090, 21204, 21318, 21432, 21546, 21660, 21774, 21888, 22002, 22116, 22230, 22344, 22458, 22572, 22686, 22800, 22914, 23028, 23142, 23256, 23370, 23484, 23598, 23712, 23826, 23940, 24054, 24168, 24282, 24396, 24510, 24624, 24738, 24852, 24966, 25080, 25194, 25308, 25422, 25536, 25650, 25764, 25878, 25992, 26106, 26220, 26334, 26448, 26562, 26676, 26790, 26904, 27018, 27132, 27246, 27360, 27474, 27588, 27702, 27816, 27930, 28044, 28158, 28272, 28386, 28500, 28614, 28728, 28842, 28956, 29070, 
0, 115, 230, 345, 460, 575, 690, 805, 920, 1035, 1150, 1265, 1380, 1495, 1610, 1725, 1840, 1955, 2070, 2185, 2300, 2415, 2530, 2645, 2760, 2875, 2990, 3105, 3220, 3335, 3450, 3565, 3680, 3795, 3910, 4025, 4140, 4255, 4370, 4485, 4600, 4715, 4830, 4945, 5060, 5175, 5290, 5405, 5520, 5635, 5750, 5865, 5980, 6095, 6210, 6325, 6440, 6555, 6670, 6785, 6900, 7015, 7130, 7245, 7360, 7475, 7590, 7705, 7820, 7935, 8050, 8165, 8280, 8395, 8510, 8625, 8740, 8855, 8970, 9085, 9200, 9315, 9430, 9545, 9660, 9775, 9890, 10005, 10120, 10235, 10350, 10465, 10580, 10695, 10810, 10925, 11040, 11155, 11270, 11385, 11500, 11615, 11730, 11845, 11960, 12075, 12190, 12305, 12420, 12535, 12650, 12765, 12880, 12995, 13110, 13225, 13340, 13455, 13570, 13685, 13800, 13915, 14030, 14145, 14260, 14375, 14490, 14605, 14720, 14835, 14950, 15065, 15180, 15295, 15410, 15525, 15640, 15755, 15870, 15985, 16100, 16215, 16330, 16445, 16560, 16675, 16790, 16905, 17020, 17135, 17250, 17365, 17480, 17595, 17710, 17825, 17940, 18055, 18170, 18285, 18400, 18515, 18630, 18745, 18860, 18975, 19090, 19205, 19320, 19435, 19550, 19665, 19780, 19895, 20010, 20125, 20240, 20355, 20470, 20585, 20700, 20815, 20930, 21045, 21160, 21275, 21390, 21505, 21620, 21735, 21850, 21965, 22080, 22195, 22310, 22425, 22540, 22655, 22770, 22885, 23000, 23115, 23230, 23345, 23460, 23575, 23690, 23805, 23920, 24035, 24150, 24265, 24380, 24495, 24610, 24725, 24840, 24955, 25070, 25185, 25300, 25415, 25530, 25645, 25760, 25875, 25990, 26105, 26220, 26335, 26450, 26565, 26680, 26795, 26910, 27025, 27140, 27255, 27370, 27485, 27600, 27715, 27830, 27945, 28060, 28175, 28290, 28405, 28520, 28635, 28750, 28865, 28980, 29095, 29210, 29325, 
0, 116, 232, 348, 464, 580, 696, 812, 928, 1044, 1160, 1276, 1392, 1508, 1624, 1740, 1856, 1972, 2088, 2204, 2320, 2436, 2552, 2668, 2784, 2900, 3016, 3132, 3248, 3364, 3480, 3596, 3712, 3828, 3944, 4060, 4176, 4292, 4408, 4524, 4640, 4756, 4872, 4988, 5104, 5220, 5336, 5452, 5568, 5684, 5800, 5916, 6032, 6148, 6264, 6380, 6496, 6612, 6728, 6844, 6960, 7076, 7192, 7308, 7424, 7540, 7656, 7772, 7888, 8004, 8120, 8236, 8352, 8468, 8584, 8700, 8816, 8932, 9048, 9164, 9280, 9396, 9512, 9628, 9744, 9860, 9976, 10092, 10208, 10324, 10440, 10556, 10672, 10788, 10904, 11020, 11136, 11252, 11368, 11484, 11600, 11716, 11832, 11948, 12064, 12180, 12296, 12412, 12528, 12644, 12760, 12876, 12992, 13108, 13224, 13340, 13456, 13572, 13688, 13804, 13920, 14036, 14152, 14268, 14384, 14500, 14616, 14732, 14848, 14964, 15080, 15196, 15312, 15428, 15544, 15660, 15776, 15892, 16008, 16124, 16240, 16356, 16472, 16588, 16704, 16820, 16936, 17052, 17168, 17284, 17400, 17516, 17632, 17748, 17864, 17980, 18096, 18212, 18328, 18444, 18560, 18676, 18792, 18908, 19024, 19140, 19256, 19372, 19488, 19604, 19720, 19836, 19952, 20068, 20184, 20300, 20416, 20532, 20648, 20764, 20880, 20996, 21112, 21228, 21344, 21460, 21576, 21692, 21808, 21924, 22040, 22156, 22272, 22388, 22504, 22620, 22736, 22852, 22968, 23084, 23200, 23316, 23432, 23548, 23664, 23780, 23896, 24012, 24128, 24244, 24360, 24476, 24592, 24708, 24824, 24940, 25056, 25172, 25288, 25404, 25520, 25636, 25752, 25868, 25984, 26100, 26216, 26332, 26448, 26564, 26680, 26796, 26912, 27028, 27144, 27260, 27376, 27492, 27608, 27724, 27840, 27956, 28072, 28188, 28304, 28420, 28536, 28652, 28768, 28884, 29000, 29116, 29232, 29348, 29464, 29580, 
0, 117, 234, 351, 468, 585, 702, 819, 936, 1053, 1170, 1287, 1404, 1521, 1638, 1755, 1872, 1989, 2106, 2223, 2340, 2457, 2574, 2691, 2808, 2925, 3042, 3159, 3276, 3393, 3510, 3627, 3744, 3861, 3978, 4095, 4212, 4329, 4446, 4563, 4680, 4797, 4914, 5031, 5148, 5265, 5382, 5499, 5616, 5733, 5850, 5967, 6084, 6201, 6318, 6435, 6552, 6669, 6786, 6903, 7020, 7137, 7254, 7371, 7488, 7605, 7722, 7839, 7956, 8073, 8190, 8307, 8424, 8541, 8658, 8775, 8892, 9009, 9126, 9243, 9360, 9477, 9594, 9711, 9828, 9945, 10062, 10179, 10296, 10413, 10530, 10647, 10764, 10881, 10998, 11115, 11232, 11349, 11466, 11583, 11700, 11817, 11934, 12051, 12168, 12285, 12402, 12519, 12636, 12753, 12870, 12987, 13104, 13221, 13338, 13455, 13572, 13689, 13806, 13923, 14040, 14157, 14274, 14391, 14508, 14625, 14742, 14859, 14976, 15093, 15210, 15327, 15444, 15561, 15678, 15795, 15912, 16029, 16146, 16263, 16380, 16497, 16614, 16731, 16848, 16965, 17082, 17199, 17316, 17433, 17550, 17667, 17784, 17901, 18018, 18135, 18252, 18369, 18486, 18603, 18720, 18837, 18954, 19071, 19188, 19305, 19422, 19539, 19656, 19773, 19890, 20007, 20124, 20241, 20358, 20475, 20592, 20709, 20826, 20943, 21060, 21177, 21294, 21411, 21528, 21645, 21762, 21879, 21996, 22113, 22230, 22347, 22464, 22581, 22698, 22815, 22932, 23049, 23166, 23283, 23400, 23517, 23634, 23751, 23868, 23985, 24102, 24219, 24336, 24453, 24570, 24687, 24804, 24921, 25038, 25155, 25272, 25389, 25506, 25623, 25740, 25857, 25974, 26091, 26208, 26325, 26442, 26559, 26676, 26793, 26910, 27027, 27144, 27261, 27378, 27495, 27612, 27729, 27846, 27963, 28080, 28197, 28314, 28431, 28548, 28665, 28782, 28899, 29016, 29133, 29250, 29367, 29484, 29601, 29718, 29835, 
0, 118, 236, 354, 472, 590, 708, 826, 944, 1062, 1180, 1298, 1416, 1534, 1652, 1770, 1888, 2006, 2124, 2242, 2360, 2478, 2596, 2714, 2832, 2950, 3068, 3186, 3304, 3422, 3540, 3658, 3776, 3894, 4012, 4130, 4248, 4366, 4484, 4602, 4720, 4838, 4956, 5074, 5192, 5310, 5428, 5546, 5664, 5782, 5900, 6018, 6136, 6254, 6372, 6490, 6608, 6726, 6844, 6962, 7080, 7198, 7316, 7434, 7552, 7670, 7788, 7906, 8024, 8142, 8260, 8378, 8496, 8614, 8732, 8850, 8968, 9086, 9204, 9322, 9440, 9558, 9676, 9794, 9912, 10030, 10148, 10266, 10384, 10502, 10620, 10738, 10856, 10974, 11092, 11210, 11328, 11446, 11564, 11682, 11800, 11918, 12036, 12154, 12272, 12390, 12508, 12626, 12744, 12862, 12980, 13098, 13216, 13334, 13452, 13570, 13688, 13806, 13924, 14042, 14160, 14278, 14396, 14514, 14632, 14750, 14868, 14986, 15104, 15222, 15340, 15458, 15576, 15694, 15812, 15930, 16048, 16166, 16284, 16402, 16520, 16638, 16756, 16874, 16992, 17110, 17228, 17346, 17464, 17582, 17700, 17818, 17936, 18054, 18172, 18290, 18408, 18526, 18644, 18762, 18880, 18998, 19116, 19234, 19352, 19470, 19588, 19706, 19824, 19942, 20060, 20178, 20296, 20414, 20532, 20650, 20768, 20886, 21004, 21122, 21240, 21358, 21476, 21594, 21712, 21830, 21948, 22066, 22184, 22302, 22420, 22538, 22656, 22774, 22892, 23010, 23128, 23246, 23364, 23482, 23600, 23718, 23836, 23954, 24072, 24190, 24308, 24426, 24544, 24662, 24780, 24898, 25016, 25134, 25252, 25370, 25488, 25606, 25724, 25842, 25960, 26078, 26196, 26314, 26432, 26550, 26668, 26786, 26904, 27022, 27140, 27258, 27376, 27494, 27612, 27730, 27848, 27966, 28084, 28202, 28320, 28438, 28556, 28674, 28792, 28910, 29028, 29146, 29264, 29382, 29500, 29618, 29736, 29854, 29972, 30090, 
0, 119, 238, 357, 476, 595, 714, 833, 952, 1071, 1190, 1309, 1428, 1547, 1666, 1785, 1904, 2023, 2142, 2261, 2380, 2499, 2618, 2737, 2856, 2975, 3094, 3213, 3332, 3451, 3570, 3689, 3808, 3927, 4046, 4165, 4284, 4403, 4522, 4641, 4760, 4879, 4998, 5117, 5236, 5355, 5474, 5593, 5712, 5831, 5950, 6069, 6188, 6307, 6426, 6545, 6664, 6783, 6902, 7021, 7140, 7259, 7378, 7497, 7616, 7735, 7854, 7973, 8092, 8211, 8330, 8449, 8568, 8687, 8806, 8925, 9044, 9163, 9282, 9401, 9520, 9639, 9758, 9877, 9996, 10115, 10234, 10353, 10472, 10591, 10710, 10829, 10948, 11067, 11186, 11305, 11424, 11543, 11662, 11781, 11900, 12019, 12138, 12257, 12376, 12495, 12614, 12733, 12852, 12971, 13090, 13209, 13328, 13447, 13566, 13685, 13804, 13923, 14042, 14161, 14280, 14399, 14518, 14637, 14756, 14875, 14994, 15113, 15232, 15351, 15470, 15589, 15708, 15827, 15946, 16065, 16184, 16303, 16422, 16541, 16660, 16779, 16898, 17017, 17136, 17255, 17374, 17493, 17612, 17731, 17850, 17969, 18088, 18207, 18326, 18445, 18564, 18683, 18802, 18921, 19040, 19159, 19278, 19397, 19516, 19635, 19754, 19873, 19992, 20111, 20230, 20349, 20468, 20587, 20706, 20825, 20944, 21063, 21182, 21301, 21420, 21539, 21658, 21777, 21896, 22015, 22134, 22253, 22372, 22491, 22610, 22729, 22848, 22967, 23086, 23205, 23324, 23443, 23562, 23681, 23800, 23919, 24038, 24157, 24276, 24395, 24514, 24633, 24752, 24871, 24990, 25109, 25228, 25347, 25466, 25585, 25704, 25823, 25942, 26061, 26180, 26299, 26418, 26537, 26656, 26775, 26894, 27013, 27132, 27251, 27370, 27489, 27608, 27727, 27846, 27965, 28084, 28203, 28322, 28441, 28560, 28679, 28798, 28917, 29036, 29155, 29274, 29393, 29512, 29631, 29750, 29869, 29988, 30107, 30226, 30345, 
0, 120, 240, 360, 480, 600, 720, 840, 960, 1080, 1200, 1320, 1440, 1560, 1680, 1800, 1920, 2040, 2160, 2280, 2400, 2520, 2640, 2760, 2880, 3000, 3120, 3240, 3360, 3480, 3600, 3720, 3840, 3960, 4080, 4200, 4320, 4440, 4560, 4680, 4800, 4920, 5040, 5160, 5280, 5400, 5520, 5640, 5760, 5880, 6000, 6120, 6240, 6360, 6480, 6600, 6720, 6840, 6960, 7080, 7200, 7320, 7440, 7560, 7680, 7800, 7920, 8040, 8160, 8280, 8400, 8520, 8640, 8760, 8880, 9000, 9120, 9240, 9360, 9480, 9600, 9720, 9840, 9960, 10080, 10200, 10320, 10440, 10560, 10680, 10800, 10920, 11040, 11160, 11280, 11400, 11520, 11640, 11760, 11880, 12000, 12120, 12240, 12360, 12480, 12600, 12720, 12840, 12960, 13080, 13200, 13320, 13440, 13560, 13680, 13800, 13920, 14040, 14160, 14280, 14400, 14520, 14640, 14760, 14880, 15000, 15120, 15240, 15360, 15480, 15600, 15720, 15840, 15960, 16080, 16200, 16320, 16440, 16560, 16680, 16800, 16920, 17040, 17160, 17280, 17400, 17520, 17640, 17760, 17880, 18000, 18120, 18240, 18360, 18480, 18600, 18720, 18840, 18960, 19080, 19200, 19320, 19440, 19560, 19680, 19800, 19920, 20040, 20160, 20280, 20400, 20520, 20640, 20760, 20880, 21000, 21120, 21240, 21360, 21480, 21600, 21720, 21840, 21960, 22080, 22200, 22320, 22440, 22560, 22680, 22800, 22920, 23040, 23160, 23280, 23400, 23520, 23640, 23760, 23880, 24000, 24120, 24240, 24360, 24480, 24600, 24720, 24840, 24960, 25080, 25200, 25320, 25440, 25560, 25680, 25800, 25920, 26040, 26160, 26280, 26400, 26520, 26640, 26760, 26880, 27000, 27120, 27240, 27360, 27480, 27600, 27720, 27840, 27960, 28080, 28200, 28320, 28440, 28560, 28680, 28800, 28920, 29040, 29160, 29280, 29400, 29520, 29640, 29760, 29880, 30000, 30120, 30240, 30360, 30480, 30600, 
0, 121, 242, 363, 484, 605, 726, 847, 968, 1089, 1210, 1331, 1452, 1573, 1694, 1815, 1936, 2057, 2178, 2299, 2420, 2541, 2662, 2783, 2904, 3025, 3146, 3267, 3388, 3509, 3630, 3751, 3872, 3993, 4114, 4235, 4356, 4477, 4598, 4719, 4840, 4961, 5082, 5203, 5324, 5445, 5566, 5687, 5808, 5929, 6050, 6171, 6292, 6413, 6534, 6655, 6776, 6897, 7018, 7139, 7260, 7381, 7502, 7623, 7744, 7865, 7986, 8107, 8228, 8349, 8470, 8591, 8712, 8833, 8954, 9075, 9196, 9317, 9438, 9559, 9680, 9801, 9922, 10043, 10164, 10285, 10406, 10527, 10648, 10769, 10890, 11011, 11132, 11253, 11374, 11495, 11616, 11737, 11858, 11979, 12100, 12221, 12342, 12463, 12584, 12705, 12826, 12947, 13068, 13189, 13310, 13431, 13552, 13673, 13794, 13915, 14036, 14157, 14278, 14399, 14520, 14641, 14762, 14883, 15004, 15125, 15246, 15367, 15488, 15609, 15730, 15851, 15972, 16093, 16214, 16335, 16456, 16577, 16698, 16819, 16940, 17061, 17182, 17303, 17424, 17545, 17666, 17787, 17908, 18029, 18150, 18271, 18392, 18513, 18634, 18755, 18876, 18997, 19118, 19239, 19360, 19481, 19602, 19723, 19844, 19965, 20086, 20207, 20328, 20449, 20570, 20691, 20812, 20933, 21054, 21175, 21296, 21417, 21538, 21659, 21780, 21901, 22022, 22143, 22264, 22385, 22506, 22627, 22748, 22869, 22990, 23111, 23232, 23353, 23474, 23595, 23716, 23837, 23958, 24079, 24200, 24321, 24442, 24563, 24684, 24805, 24926, 25047, 25168, 25289, 25410, 25531, 25652, 25773, 25894, 26015, 26136, 26257, 26378, 26499, 26620, 26741, 26862, 26983, 27104, 27225, 27346, 27467, 27588, 27709, 27830, 27951, 28072, 28193, 28314, 28435, 28556, 28677, 28798, 28919, 29040, 29161, 29282, 29403, 29524, 29645, 29766, 29887, 30008, 30129, 30250, 30371, 30492, 30613, 30734, 30855, 
0, 122, 244, 366, 488, 610, 732, 854, 976, 1098, 1220, 1342, 1464, 1586, 1708, 1830, 1952, 2074, 2196, 2318, 2440, 2562, 2684, 2806, 2928, 3050, 3172, 3294, 3416, 3538, 3660, 3782, 3904, 4026, 4148, 4270, 4392, 4514, 4636, 4758, 4880, 5002, 5124, 5246, 5368, 5490, 5612, 5734, 5856, 5978, 6100, 6222, 6344, 6466, 6588, 6710, 6832, 6954, 7076, 7198, 7320, 7442, 7564, 7686, 7808, 7930, 8052, 8174, 8296, 8418, 8540, 8662, 8784, 8906, 9028, 9150, 9272, 9394, 9516, 9638, 9760, 9882, 10004, 10126, 10248, 10370, 10492, 10614, 10736, 10858, 10980, 11102, 11224, 11346, 11468, 11590, 11712, 11834, 11956, 12078, 12200, 12322, 12444, 12566, 12688, 12810, 12932, 13054, 13176, 13298, 13420, 13542, 13664, 13786, 13908, 14030, 14152, 14274, 14396, 14518, 14640, 14762, 14884, 15006, 15128, 15250, 15372, 15494, 15616, 15738, 15860, 15982, 16104, 16226, 16348, 16470, 16592, 16714, 16836, 16958, 17080, 17202, 17324, 17446, 17568, 17690, 17812, 17934, 18056, 18178, 18300, 18422, 18544, 18666, 18788, 18910, 19032, 19154, 19276, 19398, 19520, 19642, 19764, 19886, 20008, 20130, 20252, 20374, 20496, 20618, 20740, 20862, 20984, 21106, 21228, 21350, 21472, 21594, 21716, 21838, 21960, 22082, 22204, 22326, 22448, 22570, 22692, 22814, 22936, 23058, 23180, 23302, 23424, 23546, 23668, 23790, 23912, 24034, 24156, 24278, 24400, 24522, 24644, 24766, 24888, 25010, 25132, 25254, 25376, 25498, 25620, 25742, 25864, 25986, 26108, 26230, 26352, 26474, 26596, 26718, 26840, 26962, 27084, 27206, 27328, 27450, 27572, 27694, 27816, 27938, 28060, 28182, 28304, 28426, 28548, 28670, 28792, 28914, 29036, 29158, 29280, 29402, 29524, 29646, 29768, 29890, 30012, 30134, 30256, 30378, 30500, 30622, 30744, 30866, 30988, 31110, 
0, 123, 246, 369, 492, 615, 738, 861, 984, 1107, 1230, 1353, 1476, 1599, 1722, 1845, 1968, 2091, 2214, 2337, 2460, 2583, 2706, 2829, 2952, 3075, 3198, 3321, 3444, 3567, 3690, 3813, 3936, 4059, 4182, 4305, 4428, 4551, 4674, 4797, 4920, 5043, 5166, 5289, 5412, 5535, 5658, 5781, 5904, 6027, 6150, 6273, 6396, 6519, 6642, 6765, 6888, 7011, 7134, 7257, 7380, 7503, 7626, 7749, 7872, 7995, 8118, 8241, 8364, 8487, 8610, 8733, 8856, 8979, 9102, 9225, 9348, 9471, 9594, 9717, 9840, 9963, 10086, 10209, 10332, 10455, 10578, 10701, 10824, 10947, 11070, 11193, 11316, 11439, 11562, 11685, 11808, 11931, 12054, 12177, 12300, 12423, 12546, 12669, 12792, 12915, 13038, 13161, 13284, 13407, 13530, 13653, 13776, 13899, 14022, 14145, 14268, 14391, 14514, 14637, 14760, 14883, 15006, 15129, 15252, 15375, 15498, 15621, 15744, 15867, 15990, 16113, 16236, 16359, 16482, 16605, 16728, 16851, 16974, 17097, 17220, 17343, 17466, 17589, 17712, 17835, 17958, 18081, 18204, 18327, 18450, 18573, 18696, 18819, 18942, 19065, 19188, 19311, 19434, 19557, 19680, 19803, 19926, 20049, 20172, 20295, 20418, 20541, 20664, 20787, 20910, 21033, 21156, 21279, 21402, 21525, 21648, 21771, 21894, 22017, 22140, 22263, 22386, 22509, 22632, 22755, 22878, 23001, 23124, 23247, 23370, 23493, 23616, 23739, 23862, 23985, 24108, 24231, 24354, 24477, 24600, 24723, 24846, 24969, 25092, 25215, 25338, 25461, 25584, 25707, 25830, 25953, 26076, 26199, 26322, 26445, 26568, 26691, 26814, 26937, 27060, 27183, 27306, 27429, 27552, 27675, 27798, 27921, 28044, 28167, 28290, 28413, 28536, 28659, 28782, 28905, 29028, 29151, 29274, 29397, 29520, 29643, 29766, 29889, 30012, 30135, 30258, 30381, 30504, 30627, 30750, 30873, 30996, 31119, 31242, 31365, 
0, 124, 248, 372, 496, 620, 744, 868, 992, 1116, 1240, 1364, 1488, 1612, 1736, 1860, 1984, 2108, 2232, 2356, 2480, 2604, 2728, 2852, 2976, 3100, 3224, 3348, 3472, 3596, 3720, 3844, 3968, 4092, 4216, 4340, 4464, 4588, 4712, 4836, 4960, 5084, 5208, 5332, 5456, 5580, 5704, 5828, 5952, 6076, 6200, 6324, 6448, 6572, 6696, 6820, 6944, 7068, 7192, 7316, 7440, 7564, 7688, 7812, 7936, 8060, 8184, 8308, 8432, 8556, 8680, 8804, 8928, 9052, 9176, 9300, 9424, 9548, 9672, 9796, 9920, 10044, 10168, 10292, 10416, 10540, 10664, 10788, 10912, 11036, 11160, 11284, 11408, 11532, 11656, 11780, 11904, 12028, 12152, 12276, 12400, 12524, 12648, 12772, 12896, 13020, 13144, 13268, 13392, 13516, 13640, 13764, 13888, 14012, 14136, 14260, 14384, 14508, 14632, 14756, 14880, 15004, 15128, 15252, 15376, 15500, 15624, 15748, 15872, 15996, 16120, 16244, 16368, 16492, 16616, 16740, 16864, 16988, 17112, 17236, 17360, 17484, 17608, 17732, 17856, 17980, 18104, 18228, 18352, 18476, 18600, 18724, 18848, 18972, 19096, 19220, 19344, 19468, 19592, 19716, 19840, 19964, 20088, 20212, 20336, 20460, 20584, 20708, 20832, 20956, 21080, 21204, 21328, 21452, 21576, 21700, 21824, 21948, 22072, 22196, 22320, 22444, 22568, 22692, 22816, 22940, 23064, 23188, 23312, 23436, 23560, 23684, 23808, 23932, 24056, 24180, 24304, 24428, 24552, 24676, 24800, 24924, 25048, 25172, 25296, 25420, 25544, 25668, 25792, 25916, 26040, 26164, 26288, 26412, 26536, 26660, 26784, 26908, 27032, 27156, 27280, 27404, 27528, 27652, 27776, 27900, 28024, 28148, 28272, 28396, 28520, 28644, 28768, 28892, 29016, 29140, 29264, 29388, 29512, 29636, 29760, 29884, 30008, 30132, 30256, 30380, 30504, 30628, 30752, 30876, 31000, 31124, 31248, 31372, 31496, 31620, 
0, 125, 250, 375, 500, 625, 750, 875, 1000, 1125, 1250, 1375, 1500, 1625, 1750, 1875, 2000, 2125, 2250, 2375, 2500, 2625, 2750, 2875, 3000, 3125, 3250, 3375, 3500, 3625, 3750, 3875, 4000, 4125, 4250, 4375, 4500, 4625, 4750, 4875, 5000, 5125, 5250, 5375, 5500, 5625, 5750, 5875, 6000, 6125, 6250, 6375, 6500, 6625, 6750, 6875, 7000, 7125, 7250, 7375, 7500, 7625, 7750, 7875, 8000, 8125, 8250, 8375, 8500, 8625, 8750, 8875, 9000, 9125, 9250, 9375, 9500, 9625, 9750, 9875, 10000, 10125, 10250, 10375, 10500, 10625, 10750, 10875, 11000, 11125, 11250, 11375, 11500, 11625, 11750, 11875, 12000, 12125, 12250, 12375, 12500, 12625, 12750, 12875, 13000, 13125, 13250, 13375, 13500, 13625, 13750, 13875, 14000, 14125, 14250, 14375, 14500, 14625, 14750, 14875, 15000, 15125, 15250, 15375, 15500, 15625, 15750, 15875, 16000, 16125, 16250, 16375, 16500, 16625, 16750, 16875, 17000, 17125, 17250, 17375, 17500, 17625, 17750, 17875, 18000, 18125, 18250, 18375, 18500, 18625, 18750, 18875, 19000, 19125, 19250, 19375, 19500, 19625, 19750, 19875, 20000, 20125, 20250, 20375, 20500, 20625, 20750, 20875, 21000, 21125, 21250, 21375, 21500, 21625, 21750, 21875, 22000, 22125, 22250, 22375, 22500, 22625, 22750, 22875, 23000, 23125, 23250, 23375, 23500, 23625, 23750, 23875, 24000, 24125, 24250, 24375, 24500, 24625, 24750, 24875, 25000, 25125, 25250, 25375, 25500, 25625, 25750, 25875, 26000, 26125, 26250, 26375, 26500, 26625, 26750, 26875, 27000, 27125, 27250, 27375, 27500, 27625, 27750, 27875, 28000, 28125, 28250, 28375, 28500, 28625, 28750, 28875, 29000, 29125, 29250, 29375, 29500, 29625, 29750, 29875, 30000, 30125, 30250, 30375, 30500, 30625, 30750, 30875, 31000, 31125, 31250, 31375, 31500, 31625, 31750, 31875, 
0, 126, 252, 378, 504, 630, 756, 882, 1008, 1134, 1260, 1386, 1512, 1638, 1764, 1890, 2016, 2142, 2268, 2394, 2520, 2646, 2772, 2898, 3024, 3150, 3276, 3402, 3528, 3654, 3780, 3906, 4032, 4158, 4284, 4410, 4536, 4662, 4788, 4914, 5040, 5166, 5292, 5418, 5544, 5670, 5796, 5922, 6048, 6174, 6300, 6426, 6552, 6678, 6804, 6930, 7056, 7182, 7308, 7434, 7560, 7686, 7812, 7938, 8064, 8190, 8316, 8442, 8568, 8694, 8820, 8946, 9072, 9198, 9324, 9450, 9576, 9702, 9828, 9954, 10080, 10206, 10332, 10458, 10584, 10710, 10836, 10962, 11088, 11214, 11340, 11466, 11592, 11718, 11844, 11970, 12096, 12222, 12348, 12474, 12600, 12726, 12852, 12978, 13104, 13230, 13356, 13482, 13608, 13734, 13860, 13986, 14112, 14238, 14364, 14490, 14616, 14742, 14868, 14994, 15120, 15246, 15372, 15498, 15624, 15750, 15876, 16002, 16128, 16254, 16380, 16506, 16632, 16758, 16884, 17010, 17136, 17262, 17388, 17514, 17640, 17766, 17892, 18018, 18144, 18270, 18396, 18522, 18648, 18774, 18900, 19026, 19152, 19278, 19404, 19530, 19656, 19782, 19908, 20034, 20160, 20286, 20412, 20538, 20664, 20790, 20916, 21042, 21168, 21294, 21420, 21546, 21672, 21798, 21924, 22050, 22176, 22302, 22428, 22554, 22680, 22806, 22932, 23058, 23184, 23310, 23436, 23562, 23688, 23814, 23940, 24066, 24192, 24318, 24444, 24570, 24696, 24822, 24948, 25074, 25200, 25326, 25452, 25578, 25704, 25830, 25956, 26082, 26208, 26334, 26460, 26586, 26712, 26838, 26964, 27090, 27216, 27342, 27468, 27594, 27720, 27846, 27972, 28098, 28224, 28350, 28476, 28602, 28728, 28854, 28980, 29106, 29232, 29358, 29484, 29610, 29736, 29862, 29988, 30114, 30240, 30366, 30492, 30618, 30744, 30870, 30996, 31122, 31248, 31374, 31500, 31626, 31752, 31878, 32004, 32130, 
0, 127, 254, 381, 508, 635, 762, 889, 1016, 1143, 1270, 1397, 1524, 1651, 1778, 1905, 2032, 2159, 2286, 2413, 2540, 2667, 2794, 2921, 3048, 3175, 3302, 3429, 3556, 3683, 3810, 3937, 4064, 4191, 4318, 4445, 4572, 4699, 4826, 4953, 5080, 5207, 5334, 5461, 5588, 5715, 5842, 5969, 6096, 6223, 6350, 6477, 6604, 6731, 6858, 6985, 7112, 7239, 7366, 7493, 7620, 7747, 7874, 8001, 8128, 8255, 8382, 8509, 8636, 8763, 8890, 9017, 9144, 9271, 9398, 9525, 9652, 9779, 9906, 10033, 10160, 10287, 10414, 10541, 10668, 10795, 10922, 11049, 11176, 11303, 11430, 11557, 11684, 11811, 11938, 12065, 12192, 12319, 12446, 12573, 12700, 12827, 12954, 13081, 13208, 13335, 13462, 13589, 13716, 13843, 13970, 14097, 14224, 14351, 14478, 14605, 14732, 14859, 14986, 15113, 15240, 15367, 15494, 15621, 15748, 15875, 16002, 16129, 16256, 16383, 16510, 16637, 16764, 16891, 17018, 17145, 17272, 17399, 17526, 17653, 17780, 17907, 18034, 18161, 18288, 18415, 18542, 18669, 18796, 18923, 19050, 19177, 19304, 19431, 19558, 19685, 19812, 19939, 20066, 20193, 20320, 20447, 20574, 20701, 20828, 20955, 21082, 21209, 21336, 21463, 21590, 21717, 21844, 21971, 22098, 22225, 22352, 22479, 22606, 22733, 22860, 22987, 23114, 23241, 23368, 23495, 23622, 23749, 23876, 24003, 24130, 24257, 24384, 24511, 24638, 24765, 24892, 25019, 25146, 25273, 25400, 25527, 25654, 25781, 25908, 26035, 26162, 26289, 26416, 26543, 26670, 26797, 26924, 27051, 27178, 27305, 27432, 27559, 27686, 27813, 27940, 28067, 28194, 28321, 28448, 28575, 28702, 28829, 28956, 29083, 29210, 29337, 29464, 29591, 29718, 29845, 29972, 30099, 30226, 30353, 30480, 30607, 30734, 30861, 30988, 31115, 31242, 31369, 31496, 31623, 31750, 31877, 32004, 32131, 32258, 32385, 
0, 128, 256, 384, 512, 640, 768, 896, 1024, 1152, 1280, 1408, 1536, 1664, 1792, 1920, 2048, 2176, 2304, 2432, 2560, 2688, 2816, 2944, 3072, 3200, 3328, 3456, 3584, 3712, 3840, 3968, 4096, 4224, 4352, 4480, 4608, 4736, 4864, 4992, 5120, 5248, 5376, 5504, 5632, 5760, 5888, 6016, 6144, 6272, 6400, 6528, 6656, 6784, 6912, 7040, 7168, 7296, 7424, 7552, 7680, 7808, 7936, 8064, 8192, 8320, 8448, 8576, 8704, 8832, 8960, 9088, 9216, 9344, 9472, 9600, 9728, 9856, 9984, 10112, 10240, 10368, 10496, 10624, 10752, 10880, 11008, 11136, 11264, 11392, 11520, 11648, 11776, 11904, 12032, 12160, 12288, 12416, 12544, 12672, 12800, 12928, 13056, 13184, 13312, 13440, 13568, 13696, 13824, 13952, 14080, 14208, 14336, 14464, 14592, 14720, 14848, 14976, 15104, 15232, 15360, 15488, 15616, 15744, 15872, 16000, 16128, 16256, 16384, 16512, 16640, 16768, 16896, 17024, 17152, 17280, 17408, 17536, 17664, 17792, 17920, 18048, 18176, 18304, 18432, 18560, 18688, 18816, 18944, 19072, 19200, 19328, 19456, 19584, 19712, 19840, 19968, 20096, 20224, 20352, 20480, 20608, 20736, 20864, 20992, 21120, 21248, 21376, 21504, 21632, 21760, 21888, 22016, 22144, 22272, 22400, 22528, 22656, 22784, 22912, 23040, 23168, 23296, 23424, 23552, 23680, 23808, 23936, 24064, 24192, 24320, 24448, 24576, 24704, 24832, 24960, 25088, 25216, 25344, 25472, 25600, 25728, 25856, 25984, 26112, 26240, 26368, 26496, 26624, 26752, 26880, 27008, 27136, 27264, 27392, 27520, 27648, 27776, 27904, 28032, 28160, 28288, 28416, 28544, 28672, 28800, 28928, 29056, 29184, 29312, 29440, 29568, 29696, 29824, 29952, 30080, 30208, 30336, 30464, 30592, 30720, 30848, 30976, 31104, 31232, 31360, 31488, 31616, 31744, 31872, 32000, 32128, 32256, 32384, 32512, 32640, 
0, 129, 258, 387, 516, 645, 774, 903, 1032, 1161, 1290, 1419, 1548, 1677, 1806, 1935, 2064, 2193, 2322, 2451, 2580, 2709, 2838, 2967, 3096, 3225, 3354, 3483, 3612, 3741, 3870, 3999, 4128, 4257, 4386, 4515, 4644, 4773, 4902, 5031, 5160, 5289, 5418, 5547, 5676, 5805, 5934, 6063, 6192, 6321, 6450, 6579, 6708, 6837, 6966, 7095, 7224, 7353, 7482, 7611, 7740, 7869, 7998, 8127, 8256, 8385, 8514, 8643, 8772, 8901, 9030, 9159, 9288, 9417, 9546, 9675, 9804, 9933, 10062, 10191, 10320, 10449, 10578, 10707, 10836, 10965, 11094, 11223, 11352, 11481, 11610, 11739, 11868, 11997, 12126, 12255, 12384, 12513, 12642, 12771, 12900, 13029, 13158, 13287, 13416, 13545, 13674, 13803, 13932, 14061, 14190, 14319, 14448, 14577, 14706, 14835, 14964, 15093, 15222, 15351, 15480, 15609, 15738, 15867, 15996, 16125, 16254, 16383, 16512, 16641, 16770, 16899, 17028, 17157, 17286, 17415, 17544, 17673, 17802, 17931, 18060, 18189, 18318, 18447, 18576, 18705, 18834, 18963, 19092, 19221, 19350, 19479, 19608, 19737, 19866, 19995, 20124, 20253, 20382, 20511, 20640, 20769, 20898, 21027, 21156, 21285, 21414, 21543, 21672, 21801, 21930, 22059, 22188, 22317, 22446, 22575, 22704, 22833, 22962, 23091, 23220, 23349, 23478, 23607, 23736, 23865, 23994, 24123, 24252, 24381, 24510, 24639, 24768, 24897, 25026, 25155, 25284, 25413, 25542, 25671, 25800, 25929, 26058, 26187, 26316, 26445, 26574, 26703, 26832, 26961, 27090, 27219, 27348, 27477, 27606, 27735, 27864, 27993, 28122, 28251, 28380, 28509, 28638, 28767, 28896, 29025, 29154, 29283, 29412, 29541, 29670, 29799, 29928, 30057, 30186, 30315, 30444, 30573, 30702, 30831, 30960, 31089, 31218, 31347, 31476, 31605, 31734, 31863, 31992, 32121, 32250, 32379, 32508, 32637, 32766, 32895, 
0, 130, 260, 390, 520, 650, 780, 910, 1040, 1170, 1300, 1430, 1560, 1690, 1820, 1950, 2080, 2210, 2340, 2470, 2600, 2730, 2860, 2990, 3120, 3250, 3380, 3510, 3640, 3770, 3900, 4030, 4160, 4290, 4420, 4550, 4680, 4810, 4940, 5070, 5200, 5330, 5460, 5590, 5720, 5850, 5980, 6110, 6240, 6370, 6500, 6630, 6760, 6890, 7020, 7150, 7280, 7410, 7540, 7670, 7800, 7930, 8060, 8190, 8320, 8450, 8580, 8710, 8840, 8970, 9100, 9230, 9360, 9490, 9620, 9750, 9880, 10010, 10140, 10270, 10400, 10530, 10660, 10790, 10920, 11050, 11180, 11310, 11440, 11570, 11700, 11830, 11960, 12090, 12220, 12350, 12480, 12610, 12740, 12870, 13000, 13130, 13260, 13390, 13520, 13650, 13780, 13910, 14040, 14170, 14300, 14430, 14560, 14690, 14820, 14950, 15080, 15210, 15340, 15470, 15600, 15730, 15860, 15990, 16120, 16250, 16380, 16510, 16640, 16770, 16900, 17030, 17160, 17290, 17420, 17550, 17680, 17810, 17940, 18070, 18200, 18330, 18460, 18590, 18720, 18850, 18980, 19110, 19240, 19370, 19500, 19630, 19760, 19890, 20020, 20150, 20280, 20410, 20540, 20670, 20800, 20930, 21060, 21190, 21320, 21450, 21580, 21710, 21840, 21970, 22100, 22230, 22360, 22490, 22620, 22750, 22880, 23010, 23140, 23270, 23400, 23530, 23660, 23790, 23920, 24050, 24180, 24310, 24440, 24570, 24700, 24830, 24960, 25090, 25220, 25350, 25480, 25610, 25740, 25870, 26000, 26130, 26260, 26390, 26520, 26650, 26780, 26910, 27040, 27170, 27300, 27430, 27560, 27690, 27820, 27950, 28080, 28210, 28340, 28470, 28600, 28730, 28860, 28990, 29120, 29250, 29380, 29510, 29640, 29770, 29900, 30030, 30160, 30290, 30420, 30550, 30680, 30810, 30940, 31070, 31200, 31330, 31460, 31590, 31720, 31850, 31980, 32110, 32240, 32370, 32500, 32630, 32760, 32890, 33020, 33150, 
0, 131, 262, 393, 524, 655, 786, 917, 1048, 1179, 1310, 1441, 1572, 1703, 1834, 1965, 2096, 2227, 2358, 2489, 2620, 2751, 2882, 3013, 3144, 3275, 3406, 3537, 3668, 3799, 3930, 4061, 4192, 4323, 4454, 4585, 4716, 4847, 4978, 5109, 5240, 5371, 5502, 5633, 5764, 5895, 6026, 6157, 6288, 6419, 6550, 6681, 6812, 6943, 7074, 7205, 7336, 7467, 7598, 7729, 7860, 7991, 8122, 8253, 8384, 8515, 8646, 8777, 8908, 9039, 9170, 9301, 9432, 9563, 9694, 9825, 9956, 10087, 10218, 10349, 10480, 10611, 10742, 10873, 11004, 11135, 11266, 11397, 11528, 11659, 11790, 11921, 12052, 12183, 12314, 12445, 12576, 12707, 12838, 12969, 13100, 13231, 13362, 13493, 13624, 13755, 13886, 14017, 14148, 14279, 14410, 14541, 14672, 14803, 14934, 15065, 15196, 15327, 15458, 15589, 15720, 15851, 15982, 16113, 16244, 16375, 16506, 16637, 16768, 16899, 17030, 17161, 17292, 17423, 17554, 17685, 17816, 17947, 18078, 18209, 18340, 18471, 18602, 18733, 18864, 18995, 19126, 19257, 19388, 19519, 19650, 19781, 19912, 20043, 20174, 20305, 20436, 20567, 20698, 20829, 20960, 21091, 21222, 21353, 21484, 21615, 21746, 21877, 22008, 22139, 22270, 22401, 22532, 22663, 22794, 22925, 23056, 23187, 23318, 23449, 23580, 23711, 23842, 23973, 24104, 24235, 24366, 24497, 24628, 24759, 24890, 25021, 25152, 25283, 25414, 25545, 25676, 25807, 25938, 26069, 26200, 26331, 26462, 26593, 26724, 26855, 26986, 27117, 27248, 27379, 27510, 27641, 27772, 27903, 28034, 28165, 28296, 28427, 28558, 28689, 28820, 28951, 29082, 29213, 29344, 29475, 29606, 29737, 29868, 29999, 30130, 30261, 30392, 30523, 30654, 30785, 30916, 31047, 31178, 31309, 31440, 31571, 31702, 31833, 31964, 32095, 32226, 32357, 32488, 32619, 32750, 32881, 33012, 33143, 33274, 33405, 
0, 132, 264, 396, 528, 660, 792, 924, 1056, 1188, 1320, 1452, 1584, 1716, 1848, 1980, 2112, 2244, 2376, 2508, 2640, 2772, 2904, 3036, 3168, 3300, 3432, 3564, 3696, 3828, 3960, 4092, 4224, 4356, 4488, 4620, 4752, 4884, 5016, 5148, 5280, 5412, 5544, 5676, 5808, 5940, 6072, 6204, 6336, 6468, 6600, 6732, 6864, 6996, 7128, 7260, 7392, 7524, 7656, 7788, 7920, 8052, 8184, 8316, 8448, 8580, 8712, 8844, 8976, 9108, 9240, 9372, 9504, 9636, 9768, 9900, 10032, 10164, 10296, 10428, 10560, 10692, 10824, 10956, 11088, 11220, 11352, 11484, 11616, 11748, 11880, 12012, 12144, 12276, 12408, 12540, 12672, 12804, 12936, 13068, 13200, 13332, 13464, 13596, 13728, 13860, 13992, 14124, 14256, 14388, 14520, 14652, 14784, 14916, 15048, 15180, 15312, 15444, 15576, 15708, 15840, 15972, 16104, 16236, 16368, 16500, 16632, 16764, 16896, 17028, 17160, 17292, 17424, 17556, 17688, 17820, 17952, 18084, 18216, 18348, 18480, 18612, 18744, 18876, 19008, 19140, 19272, 19404, 19536, 19668, 19800, 19932, 20064, 20196, 20328, 20460, 20592, 20724, 20856, 20988, 21120, 21252, 21384, 21516, 21648, 21780, 21912, 22044, 22176, 22308, 22440, 22572, 22704, 22836, 22968, 23100, 23232, 23364, 23496, 23628, 23760, 23892, 24024, 24156, 24288, 24420, 24552, 24684, 24816, 24948, 25080, 25212, 25344, 25476, 25608, 25740, 25872, 26004, 26136, 26268, 26400, 26532, 26664, 26796, 26928, 27060, 27192, 27324, 27456, 27588, 27720, 27852, 27984, 28116, 28248, 28380, 28512, 28644, 28776, 28908, 29040, 29172, 29304, 29436, 29568, 29700, 29832, 29964, 30096, 30228, 30360, 30492, 30624, 30756, 30888, 31020, 31152, 31284, 31416, 31548, 31680, 31812, 31944, 32076, 32208, 32340, 32472, 32604, 32736, 32868, 33000, 33132, 33264, 33396, 33528, 33660, 
0, 133, 266, 399, 532, 665, 798, 931, 1064, 1197, 1330, 1463, 1596, 1729, 1862, 1995, 2128, 2261, 2394, 2527, 2660, 2793, 2926, 3059, 3192, 3325, 3458, 3591, 3724, 3857, 3990, 4123, 4256, 4389, 4522, 4655, 4788, 4921, 5054, 5187, 5320, 5453, 5586, 5719, 5852, 5985, 6118, 6251, 6384, 6517, 6650, 6783, 6916, 7049, 7182, 7315, 7448, 7581, 7714, 7847, 7980, 8113, 8246, 8379, 8512, 8645, 8778, 8911, 9044, 9177, 9310, 9443, 9576, 9709, 9842, 9975, 10108, 10241, 10374, 10507, 10640, 10773, 10906, 11039, 11172, 11305, 11438, 11571, 11704, 11837, 11970, 12103, 12236, 12369, 12502, 12635, 12768, 12901, 13034, 13167, 13300, 13433, 13566, 13699, 13832, 13965, 14098, 14231, 14364, 14497, 14630, 14763, 14896, 15029, 15162, 15295, 15428, 15561, 15694, 15827, 15960, 16093, 16226, 16359, 16492, 16625, 16758, 16891, 17024, 17157, 17290, 17423, 17556, 17689, 17822, 17955, 18088, 18221, 18354, 18487, 18620, 18753, 18886, 19019, 19152, 19285, 19418, 19551, 19684, 19817, 19950, 20083, 20216, 20349, 20482, 20615, 20748, 20881, 21014, 21147, 21280, 21413, 21546, 21679, 21812, 21945, 22078, 22211, 22344, 22477, 22610, 22743, 22876, 23009, 23142, 23275, 23408, 23541, 23674, 23807, 23940, 24073, 24206, 24339, 24472, 24605, 24738, 24871, 25004, 25137, 25270, 25403, 25536, 25669, 25802, 25935, 26068, 26201, 26334, 26467, 26600, 26733, 26866, 26999, 27132, 27265, 27398, 27531, 27664, 27797, 27930, 28063, 28196, 28329, 28462, 28595, 28728, 28861, 28994, 29127, 29260, 29393, 29526, 29659, 29792, 29925, 30058, 30191, 30324, 30457, 30590, 30723, 30856, 30989, 31122, 31255, 31388, 31521, 31654, 31787, 31920, 32053, 32186, 32319, 32452, 32585, 32718, 32851, 32984, 33117, 33250, 33383, 33516, 33649, 33782, 33915, 
0, 134, 268, 402, 536, 670, 804, 938, 1072, 1206, 1340, 1474, 1608, 1742, 1876, 2010, 2144, 2278, 2412, 2546, 2680, 2814, 2948, 3082, 3216, 3350, 3484, 3618, 3752, 3886, 4020, 4154, 4288, 4422, 4556, 4690, 4824, 4958, 5092, 5226, 5360, 5494, 5628, 5762, 5896, 6030, 6164, 6298, 6432, 6566, 6700, 6834, 6968, 7102, 7236, 7370, 7504, 7638, 7772, 7906, 8040, 8174, 8308, 8442, 8576, 8710, 8844, 8978, 9112, 9246, 9380, 9514, 9648, 9782, 9916, 10050, 10184, 10318, 10452, 10586, 10720, 10854, 10988, 11122, 11256, 11390, 11524, 11658, 11792, 11926, 12060, 12194, 12328, 12462, 12596, 12730, 12864, 12998, 13132, 13266, 13400, 13534, 13668, 13802, 13936, 14070, 14204, 14338, 14472, 14606, 14740, 14874, 15008, 15142, 15276, 15410, 15544, 15678, 15812, 15946, 16080, 16214, 16348, 16482, 16616, 16750, 16884, 17018, 17152, 17286, 17420, 17554, 17688, 17822, 17956, 18090, 18224, 18358, 18492, 18626, 18760, 18894, 19028, 19162, 19296, 19430, 19564, 19698, 19832, 19966, 20100, 20234, 20368, 20502, 20636, 20770, 20904, 21038, 21172, 21306, 21440, 21574, 21708, 21842, 21976, 22110, 22244, 22378, 22512, 22646, 22780, 22914, 23048, 23182, 23316, 23450, 23584, 23718, 23852, 23986, 24120, 24254, 24388, 24522, 24656, 24790, 24924, 25058, 25192, 25326, 25460, 25594, 25728, 25862, 25996, 26130, 26264, 26398, 26532, 26666, 26800, 26934, 27068, 27202, 27336, 27470, 27604, 27738, 27872, 28006, 28140, 28274, 28408, 28542, 28676, 28810, 28944, 29078, 29212, 29346, 29480, 29614, 29748, 29882, 30016, 30150, 30284, 30418, 30552, 30686, 30820, 30954, 31088, 31222, 31356, 31490, 31624, 31758, 31892, 32026, 32160, 32294, 32428, 32562, 32696, 32830, 32964, 33098, 33232, 33366, 33500, 33634, 33768, 33902, 34036, 34170, 
0, 135, 270, 405, 540, 675, 810, 945, 1080, 1215, 1350, 1485, 1620, 1755, 1890, 2025, 2160, 2295, 2430, 2565, 2700, 2835, 2970, 3105, 3240, 3375, 3510, 3645, 3780, 3915, 4050, 4185, 4320, 4455, 4590, 4725, 4860, 4995, 5130, 5265, 5400, 5535, 5670, 5805, 5940, 6075, 6210, 6345, 6480, 6615, 6750, 6885, 7020, 7155, 7290, 7425, 7560, 7695, 7830, 7965, 8100, 8235, 8370, 8505, 8640, 8775, 8910, 9045, 9180, 9315, 9450, 9585, 9720, 9855, 9990, 10125, 10260, 10395, 10530, 10665, 10800, 10935, 11070, 11205, 11340, 11475, 11610, 11745, 11880, 12015, 12150, 12285, 12420, 12555, 12690, 12825, 12960, 13095, 13230, 13365, 13500, 13635, 13770, 13905, 14040, 14175, 14310, 14445, 14580, 14715, 14850, 14985, 15120, 15255, 15390, 15525, 15660, 15795, 15930, 16065, 16200, 16335, 16470, 16605, 16740, 16875, 17010, 17145, 17280, 17415, 17550, 17685, 17820, 17955, 18090, 18225, 18360, 18495, 18630, 18765, 18900, 19035, 19170, 19305, 19440, 19575, 19710, 19845, 19980, 20115, 20250, 20385, 20520, 20655, 20790, 20925, 21060, 21195, 21330, 21465, 21600, 21735, 21870, 22005, 22140, 22275, 22410, 22545, 22680, 22815, 22950, 23085, 23220, 23355, 23490, 23625, 23760, 23895, 24030, 24165, 24300, 24435, 24570, 24705, 24840, 24975, 25110, 25245, 25380, 25515, 25650, 25785, 25920, 26055, 26190, 26325, 26460, 26595, 26730, 26865, 27000, 27135, 27270, 27405, 27540, 27675, 27810, 27945, 28080, 28215, 28350, 28485, 28620, 28755, 28890, 29025, 29160, 29295, 29430, 29565, 29700, 29835, 29970, 30105, 30240, 30375, 30510, 30645, 30780, 30915, 31050, 31185, 31320, 31455, 31590, 31725, 31860, 31995, 32130, 32265, 32400, 32535, 32670, 32805, 32940, 33075, 33210, 33345, 33480, 33615, 33750, 33885, 34020, 34155, 34290, 34425, 
0, 136, 272, 408, 544, 680, 816, 952, 1088, 1224, 1360, 1496, 1632, 1768, 1904, 2040, 2176, 2312, 2448, 2584, 2720, 2856, 2992, 3128, 3264, 3400, 3536, 3672, 3808, 3944, 4080, 4216, 4352, 4488, 4624, 4760, 4896, 5032, 5168, 5304, 5440, 5576, 5712, 5848, 5984, 6120, 6256, 6392, 6528, 6664, 6800, 6936, 7072, 7208, 7344, 7480, 7616, 7752, 7888, 8024, 8160, 8296, 8432, 8568, 8704, 8840, 8976, 9112, 9248, 9384, 9520, 9656, 9792, 9928, 10064, 10200, 10336, 10472, 10608, 10744, 10880, 11016, 11152, 11288, 11424, 11560, 11696, 11832, 11968, 12104, 12240, 12376, 12512, 12648, 12784, 12920, 13056, 13192, 13328, 13464, 13600, 13736, 13872, 14008, 14144, 14280, 14416, 14552, 14688, 14824, 14960, 15096, 15232, 15368, 15504, 15640, 15776, 15912, 16048, 16184, 16320, 16456, 16592, 16728, 16864, 17000, 17136, 17272, 17408, 17544, 17680, 17816, 17952, 18088, 18224, 18360, 18496, 18632, 18768, 18904, 19040, 19176, 19312, 19448, 19584, 19720, 19856, 19992, 20128, 20264, 20400, 20536, 20672, 20808, 20944, 21080, 21216, 21352, 21488, 21624, 21760, 21896, 22032, 22168, 22304, 22440, 22576, 22712, 22848, 22984, 23120, 23256, 23392, 23528, 23664, 23800, 23936, 24072, 24208, 24344, 24480, 24616, 24752, 24888, 25024, 25160, 25296, 25432, 25568, 25704, 25840, 25976, 26112, 26248, 26384, 26520, 26656, 26792, 26928, 27064, 27200, 27336, 27472, 27608, 27744, 27880, 28016, 28152, 28288, 28424, 28560, 28696, 28832, 28968, 29104, 29240, 29376, 29512, 29648, 29784, 29920, 30056, 30192, 30328, 30464, 30600, 30736, 30872, 31008, 31144, 31280, 31416, 31552, 31688, 31824, 31960, 32096, 32232, 32368, 32504, 32640, 32776, 32912, 33048, 33184, 33320, 33456, 33592, 33728, 33864, 34000, 34136, 34272, 34408, 34544, 34680, 
0, 137, 274, 411, 548, 685, 822, 959, 1096, 1233, 1370, 1507, 1644, 1781, 1918, 2055, 2192, 2329, 2466, 2603, 2740, 2877, 3014, 3151, 3288, 3425, 3562, 3699, 3836, 3973, 4110, 4247, 4384, 4521, 4658, 4795, 4932, 5069, 5206, 5343, 5480, 5617, 5754, 5891, 6028, 6165, 6302, 6439, 6576, 6713, 6850, 6987, 7124, 7261, 7398, 7535, 7672, 7809, 7946, 8083, 8220, 8357, 8494, 8631, 8768, 8905, 9042, 9179, 9316, 9453, 9590, 9727, 9864, 10001, 10138, 10275, 10412, 10549, 10686, 10823, 10960, 11097, 11234, 11371, 11508, 11645, 11782, 11919, 12056, 12193, 12330, 12467, 12604, 12741, 12878, 13015, 13152, 13289, 13426, 13563, 13700, 13837, 13974, 14111, 14248, 14385, 14522, 14659, 14796, 14933, 15070, 15207, 15344, 15481, 15618, 15755, 15892, 16029, 16166, 16303, 16440, 16577, 16714, 16851, 16988, 17125, 17262, 17399, 17536, 17673, 17810, 17947, 18084, 18221, 18358, 18495, 18632, 18769, 18906, 19043, 19180, 19317, 19454, 19591, 19728, 19865, 20002, 20139, 20276, 20413, 20550, 20687, 20824, 20961, 21098, 21235, 21372, 21509, 21646, 21783, 21920, 22057, 22194, 22331, 22468, 22605, 22742, 22879, 23016, 23153, 23290, 23427, 23564, 23701, 23838, 23975, 24112, 24249, 24386, 24523, 24660, 24797, 24934, 25071, 25208, 25345, 25482, 25619, 25756, 25893, 26030, 26167, 26304, 26441, 26578, 26715, 26852, 26989, 27126, 27263, 27400, 27537, 27674, 27811, 27948, 28085, 28222, 28359, 28496, 28633, 28770, 28907, 29044, 29181, 29318, 29455, 29592, 29729, 29866, 30003, 30140, 30277, 30414, 30551, 30688, 30825, 30962, 31099, 31236, 31373, 31510, 31647, 31784, 31921, 32058, 32195, 32332, 32469, 32606, 32743, 32880, 33017, 33154, 33291, 33428, 33565, 33702, 33839, 33976, 34113, 34250, 34387, 34524, 34661, 34798, 34935, 
0, 138, 276, 414, 552, 690, 828, 966, 1104, 1242, 1380, 1518, 1656, 1794, 1932, 2070, 2208, 2346, 2484, 2622, 2760, 2898, 3036, 3174, 3312, 3450, 3588, 3726, 3864, 4002, 4140, 4278, 4416, 4554, 4692, 4830, 4968, 5106, 5244, 5382, 5520, 5658, 5796, 5934, 6072, 6210, 6348, 6486, 6624, 6762, 6900, 7038, 7176, 7314, 7452, 7590, 7728, 7866, 8004, 8142, 8280, 8418, 8556, 8694, 8832, 8970, 9108, 9246, 9384, 9522, 9660, 9798, 9936, 10074, 10212, 10350, 10488, 10626, 10764, 10902, 11040, 11178, 11316, 11454, 11592, 11730, 11868, 12006, 12144, 12282, 12420, 12558, 12696, 12834, 12972, 13110, 13248, 13386, 13524, 13662, 13800, 13938, 14076, 14214, 14352, 14490, 14628, 14766, 14904, 15042, 15180, 15318, 15456, 15594, 15732, 15870, 16008, 16146, 16284, 16422, 16560, 16698, 16836, 16974, 17112, 17250, 17388, 17526, 17664, 17802, 17940, 18078, 18216, 18354, 18492, 18630, 18768, 18906, 19044, 19182, 19320, 19458, 19596, 19734, 19872, 20010, 20148, 20286, 20424, 20562, 20700, 20838, 20976, 21114, 21252, 21390, 21528, 21666, 21804, 21942, 22080, 22218, 22356, 22494, 22632, 22770, 22908, 23046, 23184, 23322, 23460, 23598, 23736, 23874, 24012, 24150, 24288, 24426, 24564, 24702, 24840, 24978, 25116, 25254, 25392, 25530, 25668, 25806, 25944, 26082, 26220, 26358, 26496, 26634, 26772, 26910, 27048, 27186, 27324, 27462, 27600, 27738, 27876, 28014, 28152, 28290, 28428, 28566, 28704, 28842, 28980, 29118, 29256, 29394, 29532, 29670, 29808, 29946, 30084, 30222, 30360, 30498, 30636, 30774, 30912, 31050, 31188, 31326, 31464, 31602, 31740, 31878, 32016, 32154, 32292, 32430, 32568, 32706, 32844, 32982, 33120, 33258, 33396, 33534, 33672, 33810, 33948, 34086, 34224, 34362, 34500, 34638, 34776, 34914, 35052, 35190, 
0, 139, 278, 417, 556, 695, 834, 973, 1112, 1251, 1390, 1529, 1668, 1807, 1946, 2085, 2224, 2363, 2502, 2641, 2780, 2919, 3058, 3197, 3336, 3475, 3614, 3753, 3892, 4031, 4170, 4309, 4448, 4587, 4726, 4865, 5004, 5143, 5282, 5421, 5560, 5699, 5838, 5977, 6116, 6255, 6394, 6533, 6672, 6811, 6950, 7089, 7228, 7367, 7506, 7645, 7784, 7923, 8062, 8201, 8340, 8479, 8618, 8757, 8896, 9035, 9174, 9313, 9452, 9591, 9730, 9869, 10008, 10147, 10286, 10425, 10564, 10703, 10842, 10981, 11120, 11259, 11398, 11537, 11676, 11815, 11954, 12093, 12232, 12371, 12510, 12649, 12788, 12927, 13066, 13205, 13344, 13483, 13622, 13761, 13900, 14039, 14178, 14317, 14456, 14595, 14734, 14873, 15012, 15151, 15290, 15429, 15568, 15707, 15846, 15985, 16124, 16263, 16402, 16541, 16680, 16819, 16958, 17097, 17236, 17375, 17514, 17653, 17792, 17931, 18070, 18209, 18348, 18487, 18626, 18765, 18904, 19043, 19182, 19321, 19460, 19599, 19738, 19877, 20016, 20155, 20294, 20433, 20572, 20711, 20850, 20989, 21128, 21267, 21406, 21545, 21684, 21823, 21962, 22101, 22240, 22379, 22518, 22657, 22796, 22935, 23074, 23213, 23352, 23491, 23630, 23769, 23908, 24047, 24186, 24325, 24464, 24603, 24742, 24881, 25020, 25159, 25298, 25437, 25576, 25715, 25854, 25993, 26132, 26271, 26410, 26549, 26688, 26827, 26966, 27105, 27244, 27383, 27522, 27661, 27800, 27939, 28078, 28217, 28356, 28495, 28634, 28773, 28912, 29051, 29190, 29329, 29468, 29607, 29746, 29885, 30024, 30163, 30302, 30441, 30580, 30719, 30858, 30997, 31136, 31275, 31414, 31553, 31692, 31831, 31970, 32109, 32248, 32387, 32526, 32665, 32804, 32943, 33082, 33221, 33360, 33499, 33638, 33777, 33916, 34055, 34194, 34333, 34472, 34611, 34750, 34889, 35028, 35167, 35306, 35445, 
0, 140, 280, 420, 560, 700, 840, 980, 1120, 1260, 1400, 1540, 1680, 1820, 1960, 2100, 2240, 2380, 2520, 2660, 2800, 2940, 3080, 3220, 3360, 3500, 3640, 3780, 3920, 4060, 4200, 4340, 4480, 4620, 4760, 4900, 5040, 5180, 5320, 5460, 5600, 5740, 5880, 6020, 6160, 6300, 6440, 6580, 6720, 6860, 7000, 7140, 7280, 7420, 7560, 7700, 7840, 7980, 8120, 8260, 8400, 8540, 8680, 8820, 8960, 9100, 9240, 9380, 9520, 9660, 9800, 9940, 10080, 10220, 10360, 10500, 10640, 10780, 10920, 11060, 11200, 11340, 11480, 11620, 11760, 11900, 12040, 12180, 12320, 12460, 12600, 12740, 12880, 13020, 13160, 13300, 13440, 13580, 13720, 13860, 14000, 14140, 14280, 14420, 14560, 14700, 14840, 14980, 15120, 15260, 15400, 15540, 15680, 15820, 15960, 16100, 16240, 16380, 16520, 16660, 16800, 16940, 17080, 17220, 17360, 17500, 17640, 17780, 17920, 18060, 18200, 18340, 18480, 18620, 18760, 18900, 19040, 19180, 19320, 19460, 19600, 19740, 19880, 20020, 20160, 20300, 20440, 20580, 20720, 20860, 21000, 21140, 21280, 21420, 21560, 21700, 21840, 21980, 22120, 22260, 22400, 22540, 22680, 22820, 22960, 23100, 23240, 23380, 23520, 23660, 23800, 23940, 24080, 24220, 24360, 24500, 24640, 24780, 24920, 25060, 25200, 25340, 25480, 25620, 25760, 25900, 26040, 26180, 26320, 26460, 26600, 26740, 26880, 27020, 27160, 27300, 27440, 27580, 27720, 27860, 28000, 28140, 28280, 28420, 28560, 28700, 28840, 28980, 29120, 29260, 29400, 29540, 29680, 29820, 29960, 30100, 30240, 30380, 30520, 30660, 30800, 30940, 31080, 31220, 31360, 31500, 31640, 31780, 31920, 32060, 32200, 32340, 32480, 32620, 32760, 32900, 33040, 33180, 33320, 33460, 33600, 33740, 33880, 34020, 34160, 34300, 34440, 34580, 34720, 34860, 35000, 35140, 35280, 35420, 35560, 35700, 
0, 141, 282, 423, 564, 705, 846, 987, 1128, 1269, 1410, 1551, 1692, 1833, 1974, 2115, 2256, 2397, 2538, 2679, 2820, 2961, 3102, 3243, 3384, 3525, 3666, 3807, 3948, 4089, 4230, 4371, 4512, 4653, 4794, 4935, 5076, 5217, 5358, 5499, 5640, 5781, 5922, 6063, 6204, 6345, 6486, 6627, 6768, 6909, 7050, 7191, 7332, 7473, 7614, 7755, 7896, 8037, 8178, 8319, 8460, 8601, 8742, 8883, 9024, 9165, 9306, 9447, 9588, 9729, 9870, 10011, 10152, 10293, 10434, 10575, 10716, 10857, 10998, 11139, 11280, 11421, 11562, 11703, 11844, 11985, 12126, 12267, 12408, 12549, 12690, 12831, 12972, 13113, 13254, 13395, 13536, 13677, 13818, 13959, 14100, 14241, 14382, 14523, 14664, 14805, 14946, 15087, 15228, 15369, 15510, 15651, 15792, 15933, 16074, 16215, 16356, 16497, 16638, 16779, 16920, 17061, 17202, 17343, 17484, 17625, 17766, 17907, 18048, 18189, 18330, 18471, 18612, 18753, 18894, 19035, 19176, 19317, 19458, 19599, 19740, 19881, 20022, 20163, 20304, 20445, 20586, 20727, 20868, 21009, 21150, 21291, 21432, 21573, 21714, 21855, 21996, 22137, 22278, 22419, 22560, 22701, 22842, 22983, 23124, 23265, 23406, 23547, 23688, 23829, 23970, 24111, 24252, 24393, 24534, 24675, 24816, 24957, 25098, 25239, 25380, 25521, 25662, 25803, 25944, 26085, 26226, 26367, 26508, 26649, 26790, 26931, 27072, 27213, 27354, 27495, 27636, 27777, 27918, 28059, 28200, 28341, 28482, 28623, 28764, 28905, 29046, 29187, 29328, 29469, 29610, 29751, 29892, 30033, 30174, 30315, 30456, 30597, 30738, 30879, 31020, 31161, 31302, 31443, 31584, 31725, 31866, 32007, 32148, 32289, 32430, 32571, 32712, 32853, 32994, 33135, 33276, 33417, 33558, 33699, 33840, 33981, 34122, 34263, 34404, 34545, 34686, 34827, 34968, 35109, 35250, 35391, 35532, 35673, 35814, 35955, 
0, 142, 284, 426, 568, 710, 852, 994, 1136, 1278, 1420, 1562, 1704, 1846, 1988, 2130, 2272, 2414, 2556, 2698, 2840, 2982, 3124, 3266, 3408, 3550, 3692, 3834, 3976, 4118, 4260, 4402, 4544, 4686, 4828, 4970, 5112, 5254, 5396, 5538, 5680, 5822, 5964, 6106, 6248, 6390, 6532, 6674, 6816, 6958, 7100, 7242, 7384, 7526, 7668, 7810, 7952, 8094, 8236, 8378, 8520, 8662, 8804, 8946, 9088, 9230, 9372, 9514, 9656, 9798, 9940, 10082, 10224, 10366, 10508, 10650, 10792, 10934, 11076, 11218, 11360, 11502, 11644, 11786, 11928, 12070, 12212, 12354, 12496, 12638, 12780, 12922, 13064, 13206, 13348, 13490, 13632, 13774, 13916, 14058, 14200, 14342, 14484, 14626, 14768, 14910, 15052, 15194, 15336, 15478, 15620, 15762, 15904, 16046, 16188, 16330, 16472, 16614, 16756, 16898, 17040, 17182, 17324, 17466, 17608, 17750, 17892, 18034, 18176, 18318, 18460, 18602, 18744, 18886, 19028, 19170, 19312, 19454, 19596, 19738, 19880, 20022, 20164, 20306, 20448, 20590, 20732, 20874, 21016, 21158, 21300, 21442, 21584, 21726, 21868, 22010, 22152, 22294, 22436, 22578, 22720, 22862, 23004, 23146, 23288, 23430, 23572, 23714, 23856, 23998, 24140, 24282, 24424, 24566, 24708, 24850, 24992, 25134, 25276, 25418, 25560, 25702, 25844, 25986, 26128, 26270, 26412, 26554, 26696, 26838, 26980, 27122, 27264, 27406, 27548, 27690, 27832, 27974, 28116, 28258, 28400, 28542, 28684, 28826, 28968, 29110, 29252, 29394, 29536, 29678, 29820, 29962, 30104, 30246, 30388, 30530, 30672, 30814, 30956, 31098, 31240, 31382, 31524, 31666, 31808, 31950, 32092, 32234, 32376, 32518, 32660, 32802, 32944, 33086, 33228, 33370, 33512, 33654, 33796, 33938, 34080, 34222, 34364, 34506, 34648, 34790, 34932, 35074, 35216, 35358, 35500, 35642, 35784, 35926, 36068, 36210, 
0, 143, 286, 429, 572, 715, 858, 1001, 1144, 1287, 1430, 1573, 1716, 1859, 2002, 2145, 2288, 2431, 2574, 2717, 2860, 3003, 3146, 3289, 3432, 3575, 3718, 3861, 4004, 4147, 4290, 4433, 4576, 4719, 4862, 5005, 5148, 5291, 5434, 5577, 5720, 5863, 6006, 6149, 6292, 6435, 6578, 6721, 6864, 7007, 7150, 7293, 7436, 7579, 7722, 7865, 8008, 8151, 8294, 8437, 8580, 8723, 8866, 9009, 9152, 9295, 9438, 9581, 9724, 9867, 10010, 10153, 10296, 10439, 10582, 10725, 10868, 11011, 11154, 11297, 11440, 11583, 11726, 11869, 12012, 12155, 12298, 12441, 12584, 12727, 12870, 13013, 13156, 13299, 13442, 13585, 13728, 13871, 14014, 14157, 14300, 14443, 14586, 14729, 14872, 15015, 15158, 15301, 15444, 15587, 15730, 15873, 16016, 16159, 16302, 16445, 16588, 16731, 16874, 17017, 17160, 17303, 17446, 17589, 17732, 17875, 18018, 18161, 18304, 18447, 18590, 18733, 18876, 19019, 19162, 19305, 19448, 19591, 19734, 19877, 20020, 20163, 20306, 20449, 20592, 20735, 20878, 21021, 21164, 21307, 21450, 21593, 21736, 21879, 22022, 22165, 22308, 22451, 22594, 22737, 22880, 23023, 23166, 23309, 23452, 23595, 23738, 23881, 24024, 24167, 24310, 24453, 24596, 24739, 24882, 25025, 25168, 25311, 25454, 25597, 25740, 25883, 26026, 26169, 26312, 26455, 26598, 26741, 26884, 27027, 27170, 27313, 27456, 27599, 27742, 27885, 28028, 28171, 28314, 28457, 28600, 28743, 28886, 29029, 29172, 29315, 29458, 29601, 29744, 29887, 30030, 30173, 30316, 30459, 30602, 30745, 30888, 31031, 31174, 31317, 31460, 31603, 31746, 31889, 32032, 32175, 32318, 32461, 32604, 32747, 32890, 33033, 33176, 33319, 33462, 33605, 33748, 33891, 34034, 34177, 34320, 34463, 34606, 34749, 34892, 35035, 35178, 35321, 35464, 35607, 35750, 35893, 36036, 36179, 36322, 36465, 
0, 144, 288, 432, 576, 720, 864, 1008, 1152, 1296, 1440, 1584, 1728, 1872, 2016, 2160, 2304, 2448, 2592, 2736, 2880, 3024, 3168, 3312, 3456, 3600, 3744, 3888, 4032, 4176, 4320, 4464, 4608, 4752, 4896, 5040, 5184, 5328, 5472, 5616, 5760, 5904, 6048, 6192, 6336, 6480, 6624, 6768, 6912, 7056, 7200, 7344, 7488, 7632, 7776, 7920, 8064, 8208, 8352, 8496, 8640, 8784, 8928, 9072, 9216, 9360, 9504, 9648, 9792, 9936, 10080, 10224, 10368, 10512, 10656, 10800, 10944, 11088, 11232, 11376, 11520, 11664, 11808, 11952, 12096, 12240, 12384, 12528, 12672, 12816, 12960, 13104, 13248, 13392, 13536, 13680, 13824, 13968, 14112, 14256, 14400, 14544, 14688, 14832, 14976, 15120, 15264, 15408, 15552, 15696, 15840, 15984, 16128, 16272, 16416, 16560, 16704, 16848, 16992, 17136, 17280, 17424, 17568, 17712, 17856, 18000, 18144, 18288, 18432, 18576, 18720, 18864, 19008, 19152, 19296, 19440, 19584, 19728, 19872, 20016, 20160, 20304, 20448, 20592, 20736, 20880, 21024, 21168, 21312, 21456, 21600, 21744, 21888, 22032, 22176, 22320, 22464, 22608, 22752, 22896, 23040, 23184, 23328, 23472, 23616, 23760, 23904, 24048, 24192, 24336, 24480, 24624, 24768, 24912, 25056, 25200, 25344, 25488, 25632, 25776, 25920, 26064, 26208, 26352, 26496, 26640, 26784, 26928, 27072, 27216, 27360, 27504, 27648, 27792, 27936, 28080, 28224, 28368, 28512, 28656, 28800, 28944, 29088, 29232, 29376, 29520, 29664, 29808, 29952, 30096, 30240, 30384, 30528, 30672, 30816, 30960, 31104, 31248, 31392, 31536, 31680, 31824, 31968, 32112, 32256, 32400, 32544, 32688, 32832, 32976, 33120, 33264, 33408, 33552, 33696, 33840, 33984, 34128, 34272, 34416, 34560, 34704, 34848, 34992, 35136, 35280, 35424, 35568, 35712, 35856, 36000, 36144, 36288, 36432, 36576, 36720, 
0, 145, 290, 435, 580, 725, 870, 1015, 1160, 1305, 1450, 1595, 1740, 1885, 2030, 2175, 2320, 2465, 2610, 2755, 2900, 3045, 3190, 3335, 3480, 3625, 3770, 3915, 4060, 4205, 4350, 4495, 4640, 4785, 4930, 5075, 5220, 5365, 5510, 5655, 5800, 5945, 6090, 6235, 6380, 6525, 6670, 6815, 6960, 7105, 7250, 7395, 7540, 7685, 7830, 7975, 8120, 8265, 8410, 8555, 8700, 8845, 8990, 9135, 9280, 9425, 9570, 9715, 9860, 10005, 10150, 10295, 10440, 10585, 10730, 10875, 11020, 11165, 11310, 11455, 11600, 11745, 11890, 12035, 12180, 12325, 12470, 12615, 12760, 12905, 13050, 13195, 13340, 13485, 13630, 13775, 13920, 14065, 14210, 14355, 14500, 14645, 14790, 14935, 15080, 15225, 15370, 15515, 15660, 15805, 15950, 16095, 16240, 16385, 16530, 16675, 16820, 16965, 17110, 17255, 17400, 17545, 17690, 17835, 17980, 18125, 18270, 18415, 18560, 18705, 18850, 18995, 19140, 19285, 19430, 19575, 19720, 19865, 20010, 20155, 20300, 20445, 20590, 20735, 20880, 21025, 21170, 21315, 21460, 21605, 21750, 21895, 22040, 22185, 22330, 22475, 22620, 22765, 22910, 23055, 23200, 23345, 23490, 23635, 23780, 23925, 24070, 24215, 24360, 24505, 24650, 24795, 24940, 25085, 25230, 25375, 25520, 25665, 25810, 25955, 26100, 26245, 26390, 26535, 26680, 26825, 26970, 27115, 27260, 27405, 27550, 27695, 27840, 27985, 28130, 28275, 28420, 28565, 28710, 28855, 29000, 29145, 29290, 29435, 29580, 29725, 29870, 30015, 30160, 30305, 30450, 30595, 30740, 30885, 31030, 31175, 31320, 31465, 31610, 31755, 31900, 32045, 32190, 32335, 32480, 32625, 32770, 32915, 33060, 33205, 33350, 33495, 33640, 33785, 33930, 34075, 34220, 34365, 34510, 34655, 34800, 34945, 35090, 35235, 35380, 35525, 35670, 35815, 35960, 36105, 36250, 36395, 36540, 36685, 36830, 36975, 
0, 146, 292, 438, 584, 730, 876, 1022, 1168, 1314, 1460, 1606, 1752, 1898, 2044, 2190, 2336, 2482, 2628, 2774, 2920, 3066, 3212, 3358, 3504, 3650, 3796, 3942, 4088, 4234, 4380, 4526, 4672, 4818, 4964, 5110, 5256, 5402, 5548, 5694, 5840, 5986, 6132, 6278, 6424, 6570, 6716, 6862, 7008, 7154, 7300, 7446, 7592, 7738, 7884, 8030, 8176, 8322, 8468, 8614, 8760, 8906, 9052, 9198, 9344, 9490, 9636, 9782, 9928, 10074, 10220, 10366, 10512, 10658, 10804, 10950, 11096, 11242, 11388, 11534, 11680, 11826, 11972, 12118, 12264, 12410, 12556, 12702, 12848, 12994, 13140, 13286, 13432, 13578, 13724, 13870, 14016, 14162, 14308, 14454, 14600, 14746, 14892, 15038, 15184, 15330, 15476, 15622, 15768, 15914, 16060, 16206, 16352, 16498, 16644, 16790, 16936, 17082, 17228, 17374, 17520, 17666, 17812, 17958, 18104, 18250, 18396, 18542, 18688, 18834, 18980, 19126, 19272, 19418, 19564, 19710, 19856, 20002, 20148, 20294, 20440, 20586, 20732, 20878, 21024, 21170, 21316, 21462, 21608, 21754, 21900, 22046, 22192, 22338, 22484, 22630, 22776, 22922, 23068, 23214, 23360, 23506, 23652, 23798, 23944, 24090, 24236, 24382, 24528, 24674, 24820, 24966, 25112, 25258, 25404, 25550, 25696, 25842, 25988, 26134, 26280, 26426, 26572, 26718, 26864, 27010, 27156, 27302, 27448, 27594, 27740, 27886, 28032, 28178, 28324, 28470, 28616, 28762, 28908, 29054, 29200, 29346, 29492, 29638, 29784, 29930, 30076, 30222, 30368, 30514, 30660, 30806, 30952, 31098, 31244, 31390, 31536, 31682, 31828, 31974, 32120, 32266, 32412, 32558, 32704, 32850, 32996, 33142, 33288, 33434, 33580, 33726, 33872, 34018, 34164, 34310, 34456, 34602, 34748, 34894, 35040, 35186, 35332, 35478, 35624, 35770, 35916, 36062, 36208, 36354, 36500, 36646, 36792, 36938, 37084, 37230, 
0, 147, 294, 441, 588, 735, 882, 1029, 1176, 1323, 1470, 1617, 1764, 1911, 2058, 2205, 2352, 2499, 2646, 2793, 2940, 3087, 3234, 3381, 3528, 3675, 3822, 3969, 4116, 4263, 4410, 4557, 4704, 4851, 4998, 5145, 5292, 5439, 5586, 5733, 5880, 6027, 6174, 6321, 6468, 6615, 6762, 6909, 7056, 7203, 7350, 7497, 7644, 7791, 7938, 8085, 8232, 8379, 8526, 8673, 8820, 8967, 9114, 9261, 9408, 9555, 9702, 9849, 9996, 10143, 10290, 10437, 10584, 10731, 10878, 11025, 11172, 11319, 11466, 11613, 11760, 11907, 12054, 12201, 12348, 12495, 12642, 12789, 12936, 13083, 13230, 13377, 13524, 13671, 13818, 13965, 14112, 14259, 14406, 14553, 14700, 14847, 14994, 15141, 15288, 15435, 15582, 15729, 15876, 16023, 16170, 16317, 16464, 16611, 16758, 16905, 17052, 17199, 17346, 17493, 17640, 17787, 17934, 18081, 18228, 18375, 18522, 18669, 18816, 18963, 19110, 19257, 19404, 19551, 19698, 19845, 19992, 20139, 20286, 20433, 20580, 20727, 20874, 21021, 21168, 21315, 21462, 21609, 21756, 21903, 22050, 22197, 22344, 22491, 22638, 22785, 22932, 23079, 23226, 23373, 23520, 23667, 23814, 23961, 24108, 24255, 24402, 24549, 24696, 24843, 24990, 25137, 25284, 25431, 25578, 25725, 25872, 26019, 26166, 26313, 26460, 26607, 26754, 26901, 27048, 27195, 27342, 27489, 27636, 27783, 27930, 28077, 28224, 28371, 28518, 28665, 28812, 28959, 29106, 29253, 29400, 29547, 29694, 29841, 29988, 30135, 30282, 30429, 30576, 30723, 30870, 31017, 31164, 31311, 31458, 31605, 31752, 31899, 32046, 32193, 32340, 32487, 32634, 32781, 32928, 33075, 33222, 33369, 33516, 33663, 33810, 33957, 34104, 34251, 34398, 34545, 34692, 34839, 34986, 35133, 35280, 35427, 35574, 35721, 35868, 36015, 36162, 36309, 36456, 36603, 36750, 36897, 37044, 37191, 37338, 37485, 
0, 148, 296, 444, 592, 740, 888, 1036, 1184, 1332, 1480, 1628, 1776, 1924, 2072, 2220, 2368, 2516, 2664, 2812, 2960, 3108, 3256, 3404, 3552, 3700, 3848, 3996, 4144, 4292, 4440, 4588, 4736, 4884, 5032, 5180, 5328, 5476, 5624, 5772, 5920, 6068, 6216, 6364, 6512, 6660, 6808, 6956, 7104, 7252, 7400, 7548, 7696, 7844, 7992, 8140, 8288, 8436, 8584, 8732, 8880, 9028, 9176, 9324, 9472, 9620, 9768, 9916, 10064, 10212, 10360, 10508, 10656, 10804, 10952, 11100, 11248, 11396, 11544, 11692, 11840, 11988, 12136, 12284, 12432, 12580, 12728, 12876, 13024, 13172, 13320, 13468, 13616, 13764, 13912, 14060, 14208, 14356, 14504, 14652, 14800, 14948, 15096, 15244, 15392, 15540, 15688, 15836, 15984, 16132, 16280, 16428, 16576, 16724, 16872, 17020, 17168, 17316, 17464, 17612, 17760, 17908, 18056, 18204, 18352, 18500, 18648, 18796, 18944, 19092, 19240, 19388, 19536, 19684, 19832, 19980, 20128, 20276, 20424, 20572, 20720, 20868, 21016, 21164, 21312, 21460, 21608, 21756, 21904, 22052, 22200, 22348, 22496, 22644, 22792, 22940, 23088, 23236, 23384, 23532, 23680, 23828, 23976, 24124, 24272, 24420, 24568, 24716, 24864, 25012, 25160, 25308, 25456, 25604, 25752, 25900, 26048, 26196, 26344, 26492, 26640, 26788, 26936, 27084, 27232, 27380, 27528, 27676, 27824, 27972, 28120, 28268, 28416, 28564, 28712, 28860, 29008, 29156, 29304, 29452, 29600, 29748, 29896, 30044, 30192, 30340, 30488, 30636, 30784, 30932, 31080, 31228, 31376, 31524, 31672, 31820, 31968, 32116, 32264, 32412, 32560, 32708, 32856, 33004, 33152, 33300, 33448, 33596, 33744, 33892, 34040, 34188, 34336, 34484, 34632, 34780, 34928, 35076, 35224, 35372, 35520, 35668, 35816, 35964, 36112, 36260, 36408, 36556, 36704, 36852, 37000, 37148, 37296, 37444, 37592, 37740, 
0, 149, 298, 447, 596, 745, 894, 1043, 1192, 1341, 1490, 1639, 1788, 1937, 2086, 2235, 2384, 2533, 2682, 2831, 2980, 3129, 3278, 3427, 3576, 3725, 3874, 4023, 4172, 4321, 4470, 4619, 4768, 4917, 5066, 5215, 5364, 5513, 5662, 5811, 5960, 6109, 6258, 6407, 6556, 6705, 6854, 7003, 7152, 7301, 7450, 7599, 7748, 7897, 8046, 8195, 8344, 8493, 8642, 8791, 8940, 9089, 9238, 9387, 9536, 9685, 9834, 9983, 10132, 10281, 10430, 10579, 10728, 10877, 11026, 11175, 11324, 11473, 11622, 11771, 11920, 12069, 12218, 12367, 12516, 12665, 12814, 12963, 13112, 13261, 13410, 13559, 13708, 13857, 14006, 14155, 14304, 14453, 14602, 14751, 14900, 15049, 15198, 15347, 15496, 15645, 15794, 15943, 16092, 16241, 16390, 16539, 16688, 16837, 16986, 17135, 17284, 17433, 17582, 17731, 17880, 18029, 18178, 18327, 18476, 18625, 18774, 18923, 19072, 19221, 19370, 19519, 19668, 19817, 19966, 20115, 20264, 20413, 20562, 20711, 20860, 21009, 21158, 21307, 21456, 21605, 21754, 21903, 22052, 22201, 22350, 22499, 22648, 22797, 22946, 23095, 23244, 23393, 23542, 23691, 23840, 23989, 24138, 24287, 24436, 24585, 24734, 24883, 25032, 25181, 25330, 25479, 25628, 25777, 25926, 26075, 26224, 26373, 26522, 26671, 26820, 26969, 27118, 27267, 27416, 27565, 27714, 27863, 28012, 28161, 28310, 28459, 28608, 28757, 28906, 29055, 29204, 29353, 29502, 29651, 29800, 29949, 30098, 30247, 30396, 30545, 30694, 30843, 30992, 31141, 31290, 31439, 31588, 31737, 31886, 32035, 32184, 32333, 32482, 32631, 32780, 32929, 33078, 33227, 33376, 33525, 33674, 33823, 33972, 34121, 34270, 34419, 34568, 34717, 34866, 35015, 35164, 35313, 35462, 35611, 35760, 35909, 36058, 36207, 36356, 36505, 36654, 36803, 36952, 37101, 37250, 37399, 37548, 37697, 37846, 37995, 
0, 150, 300, 450, 600, 750, 900, 1050, 1200, 1350, 1500, 1650, 1800, 1950, 2100, 2250, 2400, 2550, 2700, 2850, 3000, 3150, 3300, 3450, 3600, 3750, 3900, 4050, 4200, 4350, 4500, 4650, 4800, 4950, 5100, 5250, 5400, 5550, 5700, 5850, 6000, 6150, 6300, 6450, 6600, 6750, 6900, 7050, 7200, 7350, 7500, 7650, 7800, 7950, 8100, 8250, 8400, 8550, 8700, 8850, 9000, 9150, 9300, 9450, 9600, 9750, 9900, 10050, 10200, 10350, 10500, 10650, 10800, 10950, 11100, 11250, 11400, 11550, 11700, 11850, 12000, 12150, 12300, 12450, 12600, 12750, 12900, 13050, 13200, 13350, 13500, 13650, 13800, 13950, 14100, 14250, 14400, 14550, 14700, 14850, 15000, 15150, 15300, 15450, 15600, 15750, 15900, 16050, 16200, 16350, 16500, 16650, 16800, 16950, 17100, 17250, 17400, 17550, 17700, 17850, 18000, 18150, 18300, 18450, 18600, 18750, 18900, 19050, 19200, 19350, 19500, 19650, 19800, 19950, 20100, 20250, 20400, 20550, 20700, 20850, 21000, 21150, 21300, 21450, 21600, 21750, 21900, 22050, 22200, 22350, 22500, 22650, 22800, 22950, 23100, 23250, 23400, 23550, 23700, 23850, 24000, 24150, 24300, 24450, 24600, 24750, 24900, 25050, 25200, 25350, 25500, 25650, 25800, 25950, 26100, 26250, 26400, 26550, 26700, 26850, 27000, 27150, 27300, 27450, 27600, 27750, 27900, 28050, 28200, 28350, 28500, 28650, 28800, 28950, 29100, 29250, 29400, 29550, 29700, 29850, 30000, 30150, 30300, 30450, 30600, 30750, 30900, 31050, 31200, 31350, 31500, 31650, 31800, 31950, 32100, 32250, 32400, 32550, 32700, 32850, 33000, 33150, 33300, 33450, 33600, 33750, 33900, 34050, 34200, 34350, 34500, 34650, 34800, 34950, 35100, 35250, 35400, 35550, 35700, 35850, 36000, 36150, 36300, 36450, 36600, 36750, 36900, 37050, 37200, 37350, 37500, 37650, 37800, 37950, 38100, 38250, 
0, 151, 302, 453, 604, 755, 906, 1057, 1208, 1359, 1510, 1661, 1812, 1963, 2114, 2265, 2416, 2567, 2718, 2869, 3020, 3171, 3322, 3473, 3624, 3775, 3926, 4077, 4228, 4379, 4530, 4681, 4832, 4983, 5134, 5285, 5436, 5587, 5738, 5889, 6040, 6191, 6342, 6493, 6644, 6795, 6946, 7097, 7248, 7399, 7550, 7701, 7852, 8003, 8154, 8305, 8456, 8607, 8758, 8909, 9060, 9211, 9362, 9513, 9664, 9815, 9966, 10117, 10268, 10419, 10570, 10721, 10872, 11023, 11174, 11325, 11476, 11627, 11778, 11929, 12080, 12231, 12382, 12533, 12684, 12835, 12986, 13137, 13288, 13439, 13590, 13741, 13892, 14043, 14194, 14345, 14496, 14647, 14798, 14949, 15100, 15251, 15402, 15553, 15704, 15855, 16006, 16157, 16308, 16459, 16610, 16761, 16912, 17063, 17214, 17365, 17516, 17667, 17818, 17969, 18120, 18271, 18422, 18573, 18724, 18875, 19026, 19177, 19328, 19479, 19630, 19781, 19932, 20083, 20234, 20385, 20536, 20687, 20838, 20989, 21140, 21291, 21442, 21593, 21744, 21895, 22046, 22197, 22348, 22499, 22650, 22801, 22952, 23103, 23254, 23405, 23556, 23707, 23858, 24009, 24160, 24311, 24462, 24613, 24764, 24915, 25066, 25217, 25368, 25519, 25670, 25821, 25972, 26123, 26274, 26425, 26576, 26727, 26878, 27029, 27180, 27331, 27482, 27633, 27784, 27935, 28086, 28237, 28388, 28539, 28690, 28841, 28992, 29143, 29294, 29445, 29596, 29747, 29898, 30049, 30200, 30351, 30502, 30653, 30804, 30955, 31106, 31257, 31408, 31559, 31710, 31861, 32012, 32163, 32314, 32465, 32616, 32767, 32918, 33069, 33220, 33371, 33522, 33673, 33824, 33975, 34126, 34277, 34428, 34579, 34730, 34881, 35032, 35183, 35334, 35485, 35636, 35787, 35938, 36089, 36240, 36391, 36542, 36693, 36844, 36995, 37146, 37297, 37448, 37599, 37750, 37901, 38052, 38203, 38354, 38505, 
0, 152, 304, 456, 608, 760, 912, 1064, 1216, 1368, 1520, 1672, 1824, 1976, 2128, 2280, 2432, 2584, 2736, 2888, 3040, 3192, 3344, 3496, 3648, 3800, 3952, 4104, 4256, 4408, 4560, 4712, 4864, 5016, 5168, 5320, 5472, 5624, 5776, 5928, 6080, 6232, 6384, 6536, 6688, 6840, 6992, 7144, 7296, 7448, 7600, 7752, 7904, 8056, 8208, 8360, 8512, 8664, 8816, 8968, 9120, 9272, 9424, 9576, 9728, 9880, 10032, 10184, 10336, 10488, 10640, 10792, 10944, 11096, 11248, 11400, 11552, 11704, 11856, 12008, 12160, 12312, 12464, 12616, 12768, 12920, 13072, 13224, 13376, 13528, 13680, 13832, 13984, 14136, 14288, 14440, 14592, 14744, 14896, 15048, 15200, 15352, 15504, 15656, 15808, 15960, 16112, 16264, 16416, 16568, 16720, 16872, 17024, 17176, 17328, 17480, 17632, 17784, 17936, 18088, 18240, 18392, 18544, 18696, 18848, 19000, 19152, 19304, 19456, 19608, 19760, 19912, 20064, 20216, 20368, 20520, 20672, 20824, 20976, 21128, 21280, 21432, 21584, 21736, 21888, 22040, 22192, 22344, 22496, 22648, 22800, 22952, 23104, 23256, 23408, 23560, 23712, 23864, 24016, 24168, 24320, 24472, 24624, 24776, 24928, 25080, 25232, 25384, 25536, 25688, 25840, 25992, 26144, 26296, 26448, 26600, 26752, 26904, 27056, 27208, 27360, 27512, 27664, 27816, 27968, 28120, 28272, 28424, 28576, 28728, 28880, 29032, 29184, 29336, 29488, 29640, 29792, 29944, 30096, 30248, 30400, 30552, 30704, 30856, 31008, 31160, 31312, 31464, 31616, 31768, 31920, 32072, 32224, 32376, 32528, 32680, 32832, 32984, 33136, 33288, 33440, 33592, 33744, 33896, 34048, 34200, 34352, 34504, 34656, 34808, 34960, 35112, 35264, 35416, 35568, 35720, 35872, 36024, 36176, 36328, 36480, 36632, 36784, 36936, 37088, 37240, 37392, 37544, 37696, 37848, 38000, 38152, 38304, 38456, 38608, 38760, 
0, 153, 306, 459, 612, 765, 918, 1071, 1224, 1377, 1530, 1683, 1836, 1989, 2142, 2295, 2448, 2601, 2754, 2907, 3060, 3213, 3366, 3519, 3672, 3825, 3978, 4131, 4284, 4437, 4590, 4743, 4896, 5049, 5202, 5355, 5508, 5661, 5814, 5967, 6120, 6273, 6426, 6579, 6732, 6885, 7038, 7191, 7344, 7497, 7650, 7803, 7956, 8109, 8262, 8415, 8568, 8721, 8874, 9027, 9180, 9333, 9486, 9639, 9792, 9945, 10098, 10251, 10404, 10557, 10710, 10863, 11016, 11169, 11322, 11475, 11628, 11781, 11934, 12087, 12240, 12393, 12546, 12699, 12852, 13005, 13158, 13311, 13464, 13617, 13770, 13923, 14076, 14229, 14382, 14535, 14688, 14841, 14994, 15147, 15300, 15453, 15606, 15759, 15912, 16065, 16218, 16371, 16524, 16677, 16830, 16983, 17136, 17289, 17442, 17595, 17748, 17901, 18054, 18207, 18360, 18513, 18666, 18819, 18972, 19125, 19278, 19431, 19584, 19737, 19890, 20043, 20196, 20349, 20502, 20655, 20808, 20961, 21114, 21267, 21420, 21573, 21726, 21879, 22032, 22185, 22338, 22491, 22644, 22797, 22950, 23103, 23256, 23409, 23562, 23715, 23868, 24021, 24174, 24327, 24480, 24633, 24786, 24939, 25092, 25245, 25398, 25551, 25704, 25857, 26010, 26163, 26316, 26469, 26622, 26775, 26928, 27081, 27234, 27387, 27540, 27693, 27846, 27999, 28152, 28305, 28458, 28611, 28764, 28917, 29070, 29223, 29376, 29529, 29682, 29835, 29988, 30141, 30294, 30447, 30600, 30753, 30906, 31059, 31212, 31365, 31518, 31671, 31824, 31977, 32130, 32283, 32436, 32589, 32742, 32895, 33048, 33201, 33354, 33507, 33660, 33813, 33966, 34119, 34272, 34425, 34578, 34731, 34884, 35037, 35190, 35343, 35496, 35649, 35802, 35955, 36108, 36261, 36414, 36567, 36720, 36873, 37026, 37179, 37332, 37485, 37638, 37791, 37944, 38097, 38250, 38403, 38556, 38709, 38862, 39015, 
0, 154, 308, 462, 616, 770, 924, 1078, 1232, 1386, 1540, 1694, 1848, 2002, 2156, 2310, 2464, 2618, 2772, 2926, 3080, 3234, 3388, 3542, 3696, 3850, 4004, 4158, 4312, 4466, 4620, 4774, 4928, 5082, 5236, 5390, 5544, 5698, 5852, 6006, 6160, 6314, 6468, 6622, 6776, 6930, 7084, 7238, 7392, 7546, 7700, 7854, 8008, 8162, 8316, 8470, 8624, 8778, 8932, 9086, 9240, 9394, 9548, 9702, 9856, 10010, 10164, 10318, 10472, 10626, 10780, 10934, 11088, 11242, 11396, 11550, 11704, 11858, 12012, 12166, 12320, 12474, 12628, 12782, 12936, 13090, 13244, 13398, 13552, 13706, 13860, 14014, 14168, 14322, 14476, 14630, 14784, 14938, 15092, 15246, 15400, 15554, 15708, 15862, 16016, 16170, 16324, 16478, 16632, 16786, 16940, 17094, 17248, 17402, 17556, 17710, 17864, 18018, 18172, 18326, 18480, 18634, 18788, 18942, 19096, 19250, 19404, 19558, 19712, 19866, 20020, 20174, 20328, 20482, 20636, 20790, 20944, 21098, 21252, 21406, 21560, 21714, 21868, 22022, 22176, 22330, 22484, 22638, 22792, 22946, 23100, 23254, 23408, 23562, 23716, 23870, 24024, 24178, 24332, 24486, 24640, 24794, 24948, 25102, 25256, 25410, 25564, 25718, 25872, 26026, 26180, 26334, 26488, 26642, 26796, 26950, 27104, 27258, 27412, 27566, 27720, 27874, 28028, 28182, 28336, 28490, 28644, 28798, 28952, 29106, 29260, 29414, 29568, 29722, 29876, 30030, 30184, 30338, 30492, 30646, 30800, 30954, 31108, 31262, 31416, 31570, 31724, 31878, 32032, 32186, 32340, 32494, 32648, 32802, 32956, 33110, 33264, 33418, 33572, 33726, 33880, 34034, 34188, 34342, 34496, 34650, 34804, 34958, 35112, 35266, 35420, 35574, 35728, 35882, 36036, 36190, 36344, 36498, 36652, 36806, 36960, 37114, 37268, 37422, 37576, 37730, 37884, 38038, 38192, 38346, 38500, 38654, 38808, 38962, 39116, 39270, 
0, 155, 310, 465, 620, 775, 930, 1085, 1240, 1395, 1550, 1705, 1860, 2015, 2170, 2325, 2480, 2635, 2790, 2945, 3100, 3255, 3410, 3565, 3720, 3875, 4030, 4185, 4340, 4495, 4650, 4805, 4960, 5115, 5270, 5425, 5580, 5735, 5890, 6045, 6200, 6355, 6510, 6665, 6820, 6975, 7130, 7285, 7440, 7595, 7750, 7905, 8060, 8215, 8370, 8525, 8680, 8835, 8990, 9145, 9300, 9455, 9610, 9765, 9920, 10075, 10230, 10385, 10540, 10695, 10850, 11005, 11160, 11315, 11470, 11625, 11780, 11935, 12090, 12245, 12400, 12555, 12710, 12865, 13020, 13175, 13330, 13485, 13640, 13795, 13950, 14105, 14260, 14415, 14570, 14725, 14880, 15035, 15190, 15345, 15500, 15655, 15810, 15965, 16120, 16275, 16430, 16585, 16740, 16895, 17050, 17205, 17360, 17515, 17670, 17825, 17980, 18135, 18290, 18445, 18600, 18755, 18910, 19065, 19220, 19375, 19530, 19685, 19840, 19995, 20150, 20305, 20460, 20615, 20770, 20925, 21080, 21235, 21390, 21545, 21700, 21855, 22010, 22165, 22320, 22475, 22630, 22785, 22940, 23095, 23250, 23405, 23560, 23715, 23870, 24025, 24180, 24335, 24490, 24645, 24800, 24955, 25110, 25265, 25420, 25575, 25730, 25885, 26040, 26195, 26350, 26505, 26660, 26815, 26970, 27125, 27280, 27435, 27590, 27745, 27900, 28055, 28210, 28365, 28520, 28675, 28830, 28985, 29140, 29295, 29450, 29605, 29760, 29915, 30070, 30225, 30380, 30535, 30690, 30845, 31000, 31155, 31310, 31465, 31620, 31775, 31930, 32085, 32240, 32395, 32550, 32705, 32860, 33015, 33170, 33325, 33480, 33635, 33790, 33945, 34100, 34255, 34410, 34565, 34720, 34875, 35030, 35185, 35340, 35495, 35650, 35805, 35960, 36115, 36270, 36425, 36580, 36735, 36890, 37045, 37200, 37355, 37510, 37665, 37820, 37975, 38130, 38285, 38440, 38595, 38750, 38905, 39060, 39215, 39370, 39525, 
0, 156, 312, 468, 624, 780, 936, 1092, 1248, 1404, 1560, 1716, 1872, 2028, 2184, 2340, 2496, 2652, 2808, 2964, 3120, 3276, 3432, 3588, 3744, 3900, 4056, 4212, 4368, 4524, 4680, 4836, 4992, 5148, 5304, 5460, 5616, 5772, 5928, 6084, 6240, 6396, 6552, 6708, 6864, 7020, 7176, 7332, 7488, 7644, 7800, 7956, 8112, 8268, 8424, 8580, 8736, 8892, 9048, 9204, 9360, 9516, 9672, 9828, 9984, 10140, 10296, 10452, 10608, 10764, 10920, 11076, 11232, 11388, 11544, 11700, 11856, 12012, 12168, 12324, 12480, 12636, 12792, 12948, 13104, 13260, 13416, 13572, 13728, 13884, 14040, 14196, 14352, 14508, 14664, 14820, 14976, 15132, 15288, 15444, 15600, 15756, 15912, 16068, 16224, 16380, 16536, 16692, 16848, 17004, 17160, 17316, 17472, 17628, 17784, 17940, 18096, 18252, 18408, 18564, 18720, 18876, 19032, 19188, 19344, 19500, 19656, 19812, 19968, 20124, 20280, 20436, 20592, 20748, 20904, 21060, 21216, 21372, 21528, 21684, 21840, 21996, 22152, 22308, 22464, 22620, 22776, 22932, 23088, 23244, 23400, 23556, 23712, 23868, 24024, 24180, 24336, 24492, 24648, 24804, 24960, 25116, 25272, 25428, 25584, 25740, 25896, 26052, 26208, 26364, 26520, 26676, 26832, 26988, 27144, 27300, 27456, 27612, 27768, 27924, 28080, 28236, 28392, 28548, 28704, 28860, 29016, 29172, 29328, 29484, 29640, 29796, 29952, 30108, 30264, 30420, 30576, 30732, 30888, 31044, 31200, 31356, 31512, 31668, 31824, 31980, 32136, 32292, 32448, 32604, 32760, 32916, 33072, 33228, 33384, 33540, 33696, 33852, 34008, 34164, 34320, 34476, 34632, 34788, 34944, 35100, 35256, 35412, 35568, 35724, 35880, 36036, 36192, 36348, 36504, 36660, 36816, 36972, 37128, 37284, 37440, 37596, 37752, 37908, 38064, 38220, 38376, 38532, 38688, 38844, 39000, 39156, 39312, 39468, 39624, 39780, 
0, 157, 314, 471, 628, 785, 942, 1099, 1256, 1413, 1570, 1727, 1884, 2041, 2198, 2355, 2512, 2669, 2826, 2983, 3140, 3297, 3454, 3611, 3768, 3925, 4082, 4239, 4396, 4553, 4710, 4867, 5024, 5181, 5338, 5495, 5652, 5809, 5966, 6123, 6280, 6437, 6594, 6751, 6908, 7065, 7222, 7379, 7536, 7693, 7850, 8007, 8164, 8321, 8478, 8635, 8792, 8949, 9106, 9263, 9420, 9577, 9734, 9891, 10048, 10205, 10362, 10519, 10676, 10833, 10990, 11147, 11304, 11461, 11618, 11775, 11932, 12089, 12246, 12403, 12560, 12717, 12874, 13031, 13188, 13345, 13502, 13659, 13816, 13973, 14130, 14287, 14444, 14601, 14758, 14915, 15072, 15229, 15386, 15543, 15700, 15857, 16014, 16171, 16328, 16485, 16642, 16799, 16956, 17113, 17270, 17427, 17584, 17741, 17898, 18055, 18212, 18369, 18526, 18683, 18840, 18997, 19154, 19311, 19468, 19625, 19782, 19939, 20096, 20253, 20410, 20567, 20724, 20881, 21038, 21195, 21352, 21509, 21666, 21823, 21980, 22137, 22294, 22451, 22608, 22765, 22922, 23079, 23236, 23393, 23550, 23707, 23864, 24021, 24178, 24335, 24492, 24649, 24806, 24963, 25120, 25277, 25434, 25591, 25748, 25905, 26062, 26219, 26376, 26533, 26690, 26847, 27004, 27161, 27318, 27475, 27632, 27789, 27946, 28103, 28260, 28417, 28574, 28731, 28888, 29045, 29202, 29359, 29516, 29673, 29830, 29987, 30144, 30301, 30458, 30615, 30772, 30929, 31086, 31243, 31400, 31557, 31714, 31871, 32028, 32185, 32342, 32499, 32656, 32813, 32970, 33127, 33284, 33441, 33598, 33755, 33912, 34069, 34226, 34383, 34540, 34697, 34854, 35011, 35168, 35325, 35482, 35639, 35796, 35953, 36110, 36267, 36424, 36581, 36738, 36895, 37052, 37209, 37366, 37523, 37680, 37837, 37994, 38151, 38308, 38465, 38622, 38779, 38936, 39093, 39250, 39407, 39564, 39721, 39878, 40035, 
0, 158, 316, 474, 632, 790, 948, 1106, 1264, 1422, 1580, 1738, 1896, 2054, 2212, 2370, 2528, 2686, 2844, 3002, 3160, 3318, 3476, 3634, 3792, 3950, 4108, 4266, 4424, 4582, 4740, 4898, 5056, 5214, 5372, 5530, 5688, 5846, 6004, 6162, 6320, 6478, 6636, 6794, 6952, 7110, 7268, 7426, 7584, 7742, 7900, 8058, 8216, 8374, 8532, 8690, 8848, 9006, 9164, 9322, 9480, 9638, 9796, 9954, 10112, 10270, 10428, 10586, 10744, 10902, 11060, 11218, 11376, 11534, 11692, 11850, 12008, 12166, 12324, 12482, 12640, 12798, 12956, 13114, 13272, 13430, 13588, 13746, 13904, 14062, 14220, 14378, 14536, 14694, 14852, 15010, 15168, 15326, 15484, 15642, 15800, 15958, 16116, 16274, 16432, 16590, 16748, 16906, 17064, 17222, 17380, 17538, 17696, 17854, 18012, 18170, 18328, 18486, 18644, 18802, 18960, 19118, 19276, 19434, 19592, 19750, 19908, 20066, 20224, 20382, 20540, 20698, 20856, 21014, 21172, 21330, 21488, 21646, 21804, 21962, 22120, 22278, 22436, 22594, 22752, 22910, 23068, 23226, 23384, 23542, 23700, 23858, 24016, 24174, 24332, 24490, 24648, 24806, 24964, 25122, 25280, 25438, 25596, 25754, 25912, 26070, 26228, 26386, 26544, 26702, 26860, 27018, 27176, 27334, 27492, 27650, 27808, 27966, 28124, 28282, 28440, 28598, 28756, 28914, 29072, 29230, 29388, 29546, 29704, 29862, 30020, 30178, 30336, 30494, 30652, 30810, 30968, 31126, 31284, 31442, 31600, 31758, 31916, 32074, 32232, 32390, 32548, 32706, 32864, 33022, 33180, 33338, 33496, 33654, 33812, 33970, 34128, 34286, 34444, 34602, 34760, 34918, 35076, 35234, 35392, 35550, 35708, 35866, 36024, 36182, 36340, 36498, 36656, 36814, 36972, 37130, 37288, 37446, 37604, 37762, 37920, 38078, 38236, 38394, 38552, 38710, 38868, 39026, 39184, 39342, 39500, 39658, 39816, 39974, 40132, 40290, 
0, 159, 318, 477, 636, 795, 954, 1113, 1272, 1431, 1590, 1749, 1908, 2067, 2226, 2385, 2544, 2703, 2862, 3021, 3180, 3339, 3498, 3657, 3816, 3975, 4134, 4293, 4452, 4611, 4770, 4929, 5088, 5247, 5406, 5565, 5724, 5883, 6042, 6201, 6360, 6519, 6678, 6837, 6996, 7155, 7314, 7473, 7632, 7791, 7950, 8109, 8268, 8427, 8586, 8745, 8904, 9063, 9222, 9381, 9540, 9699, 9858, 10017, 10176, 10335, 10494, 10653, 10812, 10971, 11130, 11289, 11448, 11607, 11766, 11925, 12084, 12243, 12402, 12561, 12720, 12879, 13038, 13197, 13356, 13515, 13674, 13833, 13992, 14151, 14310, 14469, 14628, 14787, 14946, 15105, 15264, 15423, 15582, 15741, 15900, 16059, 16218, 16377, 16536, 16695, 16854, 17013, 17172, 17331, 17490, 17649, 17808, 17967, 18126, 18285, 18444, 18603, 18762, 18921, 19080, 19239, 19398, 19557, 19716, 19875, 20034, 20193, 20352, 20511, 20670, 20829, 20988, 21147, 21306, 21465, 21624, 21783, 21942, 22101, 22260, 22419, 22578, 22737, 22896, 23055, 23214, 23373, 23532, 23691, 23850, 24009, 24168, 24327, 24486, 24645, 24804, 24963, 25122, 25281, 25440, 25599, 25758, 25917, 26076, 26235, 26394, 26553, 26712, 26871, 27030, 27189, 27348, 27507, 27666, 27825, 27984, 28143, 28302, 28461, 28620, 28779, 28938, 29097, 29256, 29415, 29574, 29733, 29892, 30051, 30210, 30369, 30528, 30687, 30846, 31005, 31164, 31323, 31482, 31641, 31800, 31959, 32118, 32277, 32436, 32595, 32754, 32913, 33072, 33231, 33390, 33549, 33708, 33867, 34026, 34185, 34344, 34503, 34662, 34821, 34980, 35139, 35298, 35457, 35616, 35775, 35934, 36093, 36252, 36411, 36570, 36729, 36888, 37047, 37206, 37365, 37524, 37683, 37842, 38001, 38160, 38319, 38478, 38637, 38796, 38955, 39114, 39273, 39432, 39591, 39750, 39909, 40068, 40227, 40386, 40545, 
0, 160, 320, 480, 640, 800, 960, 1120, 1280, 1440, 1600, 1760, 1920, 2080, 2240, 2400, 2560, 2720, 2880, 3040, 3200, 3360, 3520, 3680, 3840, 4000, 4160, 4320, 4480, 4640, 4800, 4960, 5120, 5280, 5440, 5600, 5760, 5920, 6080, 6240, 6400, 6560, 6720, 6880, 7040, 7200, 7360, 7520, 7680, 7840, 8000, 8160, 8320, 8480, 8640, 8800, 8960, 9120, 9280, 9440, 9600, 9760, 9920, 10080, 10240, 10400, 10560, 10720, 10880, 11040, 11200, 11360, 11520, 11680, 11840, 12000, 12160, 12320, 12480, 12640, 12800, 12960, 13120, 13280, 13440, 13600, 13760, 13920, 14080, 14240, 14400, 14560, 14720, 14880, 15040, 15200, 15360, 15520, 15680, 15840, 16000, 16160, 16320, 16480, 16640, 16800, 16960, 17120, 17280, 17440, 17600, 17760, 17920, 18080, 18240, 18400, 18560, 18720, 18880, 19040, 19200, 19360, 19520, 19680, 19840, 20000, 20160, 20320, 20480, 20640, 20800, 20960, 21120, 21280, 21440, 21600, 21760, 21920, 22080, 22240, 22400, 22560, 22720, 22880, 23040, 23200, 23360, 23520, 23680, 23840, 24000, 24160, 24320, 24480, 24640, 24800, 24960, 25120, 25280, 25440, 25600, 25760, 25920, 26080, 26240, 26400, 26560, 26720, 26880, 27040, 27200, 27360, 27520, 27680, 27840, 28000, 28160, 28320, 28480, 28640, 28800, 28960, 29120, 29280, 29440, 29600, 29760, 29920, 30080, 30240, 30400, 30560, 30720, 30880, 31040, 31200, 31360, 31520, 31680, 31840, 32000, 32160, 32320, 32480, 32640, 32800, 32960, 33120, 33280, 33440, 33600, 33760, 33920, 34080, 34240, 34400, 34560, 34720, 34880, 35040, 35200, 35360, 35520, 35680, 35840, 36000, 36160, 36320, 36480, 36640, 36800, 36960, 37120, 37280, 37440, 37600, 37760, 37920, 38080, 38240, 38400, 38560, 38720, 38880, 39040, 39200, 39360, 39520, 39680, 39840, 40000, 40160, 40320, 40480, 40640, 40800, 
0, 161, 322, 483, 644, 805, 966, 1127, 1288, 1449, 1610, 1771, 1932, 2093, 2254, 2415, 2576, 2737, 2898, 3059, 3220, 3381, 3542, 3703, 3864, 4025, 4186, 4347, 4508, 4669, 4830, 4991, 5152, 5313, 5474, 5635, 5796, 5957, 6118, 6279, 6440, 6601, 6762, 6923, 7084, 7245, 7406, 7567, 7728, 7889, 8050, 8211, 8372, 8533, 8694, 8855, 9016, 9177, 9338, 9499, 9660, 9821, 9982, 10143, 10304, 10465, 10626, 10787, 10948, 11109, 11270, 11431, 11592, 11753, 11914, 12075, 12236, 12397, 12558, 12719, 12880, 13041, 13202, 13363, 13524, 13685, 13846, 14007, 14168, 14329, 14490, 14651, 14812, 14973, 15134, 15295, 15456, 15617, 15778, 15939, 16100, 16261, 16422, 16583, 16744, 16905, 17066, 17227, 17388, 17549, 17710, 17871, 18032, 18193, 18354, 18515, 18676, 18837, 18998, 19159, 19320, 19481, 19642, 19803, 19964, 20125, 20286, 20447, 20608, 20769, 20930, 21091, 21252, 21413, 21574, 21735, 21896, 22057, 22218, 22379, 22540, 22701, 22862, 23023, 23184, 23345, 23506, 23667, 23828, 23989, 24150, 24311, 24472, 24633, 24794, 24955, 25116, 25277, 25438, 25599, 25760, 25921, 26082, 26243, 26404, 26565, 26726, 26887, 27048, 27209, 27370, 27531, 27692, 27853, 28014, 28175, 28336, 28497, 28658, 28819, 28980, 29141, 29302, 29463, 29624, 29785, 29946, 30107, 30268, 30429, 30590, 30751, 30912, 31073, 31234, 31395, 31556, 31717, 31878, 32039, 32200, 32361, 32522, 32683, 32844, 33005, 33166, 33327, 33488, 33649, 33810, 33971, 34132, 34293, 34454, 34615, 34776, 34937, 35098, 35259, 35420, 35581, 35742, 35903, 36064, 36225, 36386, 36547, 36708, 36869, 37030, 37191, 37352, 37513, 37674, 37835, 37996, 38157, 38318, 38479, 38640, 38801, 38962, 39123, 39284, 39445, 39606, 39767, 39928, 40089, 40250, 40411, 40572, 40733, 40894, 41055, 
0, 162, 324, 486, 648, 810, 972, 1134, 1296, 1458, 1620, 1782, 1944, 2106, 2268, 2430, 2592, 2754, 2916, 3078, 3240, 3402, 3564, 3726, 3888, 4050, 4212, 4374, 4536, 4698, 4860, 5022, 5184, 5346, 5508, 5670, 5832, 5994, 6156, 6318, 6480, 6642, 6804, 6966, 7128, 7290, 7452, 7614, 7776, 7938, 8100, 8262, 8424, 8586, 8748, 8910, 9072, 9234, 9396, 9558, 9720, 9882, 10044, 10206, 10368, 10530, 10692, 10854, 11016, 11178, 11340, 11502, 11664, 11826, 11988, 12150, 12312, 12474, 12636, 12798, 12960, 13122, 13284, 13446, 13608, 13770, 13932, 14094, 14256, 14418, 14580, 14742, 14904, 15066, 15228, 15390, 15552, 15714, 15876, 16038, 16200, 16362, 16524, 16686, 16848, 17010, 17172, 17334, 17496, 17658, 17820, 17982, 18144, 18306, 18468, 18630, 18792, 18954, 19116, 19278, 19440, 19602, 19764, 19926, 20088, 20250, 20412, 20574, 20736, 20898, 21060, 21222, 21384, 21546, 21708, 21870, 22032, 22194, 22356, 22518, 22680, 22842, 23004, 23166, 23328, 23490, 23652, 23814, 23976, 24138, 24300, 24462, 24624, 24786, 24948, 25110, 25272, 25434, 25596, 25758, 25920, 26082, 26244, 26406, 26568, 26730, 26892, 27054, 27216, 27378, 27540, 27702, 27864, 28026, 28188, 28350, 28512, 28674, 28836, 28998, 29160, 29322, 29484, 29646, 29808, 29970, 30132, 30294, 30456, 30618, 30780, 30942, 31104, 31266, 31428, 31590, 31752, 31914, 32076, 32238, 32400, 32562, 32724, 32886, 33048, 33210, 33372, 33534, 33696, 33858, 34020, 34182, 34344, 34506, 34668, 34830, 34992, 35154, 35316, 35478, 35640, 35802, 35964, 36126, 36288, 36450, 36612, 36774, 36936, 37098, 37260, 37422, 37584, 37746, 37908, 38070, 38232, 38394, 38556, 38718, 38880, 39042, 39204, 39366, 39528, 39690, 39852, 40014, 40176, 40338, 40500, 40662, 40824, 40986, 41148, 41310, 
0, 163, 326, 489, 652, 815, 978, 1141, 1304, 1467, 1630, 1793, 1956, 2119, 2282, 2445, 2608, 2771, 2934, 3097, 3260, 3423, 3586, 3749, 3912, 4075, 4238, 4401, 4564, 4727, 4890, 5053, 5216, 5379, 5542, 5705, 5868, 6031, 6194, 6357, 6520, 6683, 6846, 7009, 7172, 7335, 7498, 7661, 7824, 7987, 8150, 8313, 8476, 8639, 8802, 8965, 9128, 9291, 9454, 9617, 9780, 9943, 10106, 10269, 10432, 10595, 10758, 10921, 11084, 11247, 11410, 11573, 11736, 11899, 12062, 12225, 12388, 12551, 12714, 12877, 13040, 13203, 13366, 13529, 13692, 13855, 14018, 14181, 14344, 14507, 14670, 14833, 14996, 15159, 15322, 15485, 15648, 15811, 15974, 16137, 16300, 16463, 16626, 16789, 16952, 17115, 17278, 17441, 17604, 17767, 17930, 18093, 18256, 18419, 18582, 18745, 18908, 19071, 19234, 19397, 19560, 19723, 19886, 20049, 20212, 20375, 20538, 20701, 20864, 21027, 21190, 21353, 21516, 21679, 21842, 22005, 22168, 22331, 22494, 22657, 22820, 22983, 23146, 23309, 23472, 23635, 23798, 23961, 24124, 24287, 24450, 24613, 24776, 24939, 25102, 25265, 25428, 25591, 25754, 25917, 26080, 26243, 26406, 26569, 26732, 26895, 27058, 27221, 27384, 27547, 27710, 27873, 28036, 28199, 28362, 28525, 28688, 28851, 29014, 29177, 29340, 29503, 29666, 29829, 29992, 30155, 30318, 30481, 30644, 30807, 30970, 31133, 31296, 31459, 31622, 31785, 31948, 32111, 32274, 32437, 32600, 32763, 32926, 33089, 33252, 33415, 33578, 33741, 33904, 34067, 34230, 34393, 34556, 34719, 34882, 35045, 35208, 35371, 35534, 35697, 35860, 36023, 36186, 36349, 36512, 36675, 36838, 37001, 37164, 37327, 37490, 37653, 37816, 37979, 38142, 38305, 38468, 38631, 38794, 38957, 39120, 39283, 39446, 39609, 39772, 39935, 40098, 40261, 40424, 40587, 40750, 40913, 41076, 41239, 41402, 41565, 
0, 164, 328, 492, 656, 820, 984, 1148, 1312, 1476, 1640, 1804, 1968, 2132, 2296, 2460, 2624, 2788, 2952, 3116, 3280, 3444, 3608, 3772, 3936, 4100, 4264, 4428, 4592, 4756, 4920, 5084, 5248, 5412, 5576, 5740, 5904, 6068, 6232, 6396, 6560, 6724, 6888, 7052, 7216, 7380, 7544, 7708, 7872, 8036, 8200, 8364, 8528, 8692, 8856, 9020, 9184, 9348, 9512, 9676, 9840, 10004, 10168, 10332, 10496, 10660, 10824, 10988, 11152, 11316, 11480, 11644, 11808, 11972, 12136, 12300, 12464, 12628, 12792, 12956, 13120, 13284, 13448, 13612, 13776, 13940, 14104, 14268, 14432, 14596, 14760, 14924, 15088, 15252, 15416, 15580, 15744, 15908, 16072, 16236, 16400, 16564, 16728, 16892, 17056, 17220, 17384, 17548, 17712, 17876, 18040, 18204, 18368, 18532, 18696, 18860, 19024, 19188, 19352, 19516, 19680, 19844, 20008, 20172, 20336, 20500, 20664, 20828, 20992, 21156, 21320, 21484, 21648, 21812, 21976, 22140, 22304, 22468, 22632, 22796, 22960, 23124, 23288, 23452, 23616, 23780, 23944, 24108, 24272, 24436, 24600, 24764, 24928, 25092, 25256, 25420, 25584, 25748, 25912, 26076, 26240, 26404, 26568, 26732, 26896, 27060, 27224, 27388, 27552, 27716, 27880, 28044, 28208, 28372, 28536, 28700, 28864, 29028, 29192, 29356, 29520, 29684, 29848, 30012, 30176, 30340, 30504, 30668, 30832, 30996, 31160, 31324, 31488, 31652, 31816, 31980, 32144, 32308, 32472, 32636, 32800, 32964, 33128, 33292, 33456, 33620, 33784, 33948, 34112, 34276, 34440, 34604, 34768, 34932, 35096, 35260, 35424, 35588, 35752, 35916, 36080, 36244, 36408, 36572, 36736, 36900, 37064, 37228, 37392, 37556, 37720, 37884, 38048, 38212, 38376, 38540, 38704, 38868, 39032, 39196, 39360, 39524, 39688, 39852, 40016, 40180, 40344, 40508, 40672, 40836, 41000, 41164, 41328, 41492, 41656, 41820, 
0, 165, 330, 495, 660, 825, 990, 1155, 1320, 1485, 1650, 1815, 1980, 2145, 2310, 2475, 2640, 2805, 2970, 3135, 3300, 3465, 3630, 3795, 3960, 4125, 4290, 4455, 4620, 4785, 4950, 5115, 5280, 5445, 5610, 5775, 5940, 6105, 6270, 6435, 6600, 6765, 6930, 7095, 7260, 7425, 7590, 7755, 7920, 8085, 8250, 8415, 8580, 8745, 8910, 9075, 9240, 9405, 9570, 9735, 9900, 10065, 10230, 10395, 10560, 10725, 10890, 11055, 11220, 11385, 11550, 11715, 11880, 12045, 12210, 12375, 12540, 12705, 12870, 13035, 13200, 13365, 13530, 13695, 13860, 14025, 14190, 14355, 14520, 14685, 14850, 15015, 15180, 15345, 15510, 15675, 15840, 16005, 16170, 16335, 16500, 16665, 16830, 16995, 17160, 17325, 17490, 17655, 17820, 17985, 18150, 18315, 18480, 18645, 18810, 18975, 19140, 19305, 19470, 19635, 19800, 19965, 20130, 20295, 20460, 20625, 20790, 20955, 21120, 21285, 21450, 21615, 21780, 21945, 22110, 22275, 22440, 22605, 22770, 22935, 23100, 23265, 23430, 23595, 23760, 23925, 24090, 24255, 24420, 24585, 24750, 24915, 25080, 25245, 25410, 25575, 25740, 25905, 26070, 26235, 26400, 26565, 26730, 26895, 27060, 27225, 27390, 27555, 27720, 27885, 28050, 28215, 28380, 28545, 28710, 28875, 29040, 29205, 29370, 29535, 29700, 29865, 30030, 30195, 30360, 30525, 30690, 30855, 31020, 31185, 31350, 31515, 31680, 31845, 32010, 32175, 32340, 32505, 32670, 32835, 33000, 33165, 33330, 33495, 33660, 33825, 33990, 34155, 34320, 34485, 34650, 34815, 34980, 35145, 35310, 35475, 35640, 35805, 35970, 36135, 36300, 36465, 36630, 36795, 36960, 37125, 37290, 37455, 37620, 37785, 37950, 38115, 38280, 38445, 38610, 38775, 38940, 39105, 39270, 39435, 39600, 39765, 39930, 40095, 40260, 40425, 40590, 40755, 40920, 41085, 41250, 41415, 41580, 41745, 41910, 42075, 
0, 166, 332, 498, 664, 830, 996, 1162, 1328, 1494, 1660, 1826, 1992, 2158, 2324, 2490, 2656, 2822, 2988, 3154, 3320, 3486, 3652, 3818, 3984, 4150, 4316, 4482, 4648, 4814, 4980, 5146, 5312, 5478, 5644, 5810, 5976, 6142, 6308, 6474, 6640, 6806, 6972, 7138, 7304, 7470, 7636, 7802, 7968, 8134, 8300, 8466, 8632, 8798, 8964, 9130, 9296, 9462, 9628, 9794, 9960, 10126, 10292, 10458, 10624, 10790, 10956, 11122, 11288, 11454, 11620, 11786, 11952, 12118, 12284, 12450, 12616, 12782, 12948, 13114, 13280, 13446, 13612, 13778, 13944, 14110, 14276, 14442, 14608, 14774, 14940, 15106, 15272, 15438, 15604, 15770, 15936, 16102, 16268, 16434, 16600, 16766, 16932, 17098, 17264, 17430, 17596, 17762, 17928, 18094, 18260, 18426, 18592, 18758, 18924, 19090, 19256, 19422, 19588, 19754, 19920, 20086, 20252, 20418, 20584, 20750, 20916, 21082, 21248, 21414, 21580, 21746, 21912, 22078, 22244, 22410, 22576, 22742, 22908, 23074, 23240, 23406, 23572, 23738, 23904, 24070, 24236, 24402, 24568, 24734, 24900, 25066, 25232, 25398, 25564, 25730, 25896, 26062, 26228, 26394, 26560, 26726, 26892, 27058, 27224, 27390, 27556, 27722, 27888, 28054, 28220, 28386, 28552, 28718, 28884, 29050, 29216, 29382, 29548, 29714, 29880, 30046, 30212, 30378, 30544, 30710, 30876, 31042, 31208, 31374, 31540, 31706, 31872, 32038, 32204, 32370, 32536, 32702, 32868, 33034, 33200, 33366, 33532, 33698, 33864, 34030, 34196, 34362, 34528, 34694, 34860, 35026, 35192, 35358, 35524, 35690, 35856, 36022, 36188, 36354, 36520, 36686, 36852, 37018, 37184, 37350, 37516, 37682, 37848, 38014, 38180, 38346, 38512, 38678, 38844, 39010, 39176, 39342, 39508, 39674, 39840, 40006, 40172, 40338, 40504, 40670, 40836, 41002, 41168, 41334, 41500, 41666, 41832, 41998, 42164, 42330, 
0, 167, 334, 501, 668, 835, 1002, 1169, 1336, 1503, 1670, 1837, 2004, 2171, 2338, 2505, 2672, 2839, 3006, 3173, 3340, 3507, 3674, 3841, 4008, 4175, 4342, 4509, 4676, 4843, 5010, 5177, 5344, 5511, 5678, 5845, 6012, 6179, 6346, 6513, 6680, 6847, 7014, 7181, 7348, 7515, 7682, 7849, 8016, 8183, 8350, 8517, 8684, 8851, 9018, 9185, 9352, 9519, 9686, 9853, 10020, 10187, 10354, 10521, 10688, 10855, 11022, 11189, 11356, 11523, 11690, 11857, 12024, 12191, 12358, 12525, 12692, 12859, 13026, 13193, 13360, 13527, 13694, 13861, 14028, 14195, 14362, 14529, 14696, 14863, 15030, 15197, 15364, 15531, 15698, 15865, 16032, 16199, 16366, 16533, 16700, 16867, 17034, 17201, 17368, 17535, 17702, 17869, 18036, 18203, 18370, 18537, 18704, 18871, 19038, 19205, 19372, 19539, 19706, 19873, 20040, 20207, 20374, 20541, 20708, 20875, 21042, 21209, 21376, 21543, 21710, 21877, 22044, 22211, 22378, 22545, 22712, 22879, 23046, 23213, 23380, 23547, 23714, 23881, 24048, 24215, 24382, 24549, 24716, 24883, 25050, 25217, 25384, 25551, 25718, 25885, 26052, 26219, 26386, 26553, 26720, 26887, 27054, 27221, 27388, 27555, 27722, 27889, 28056, 28223, 28390, 28557, 28724, 28891, 29058, 29225, 29392, 29559, 29726, 29893, 30060, 30227, 30394, 30561, 30728, 30895, 31062, 31229, 31396, 31563, 31730, 31897, 32064, 32231, 32398, 32565, 32732, 32899, 33066, 33233, 33400, 33567, 33734, 33901, 34068, 34235, 34402, 34569, 34736, 34903, 35070, 35237, 35404, 35571, 35738, 35905, 36072, 36239, 36406, 36573, 36740, 36907, 37074, 37241, 37408, 37575, 37742, 37909, 38076, 38243, 38410, 38577, 38744, 38911, 39078, 39245, 39412, 39579, 39746, 39913, 40080, 40247, 40414, 40581, 40748, 40915, 41082, 41249, 41416, 41583, 41750, 41917, 42084, 42251, 42418, 42585, 
0, 168, 336, 504, 672, 840, 1008, 1176, 1344, 1512, 1680, 1848, 2016, 2184, 2352, 2520, 2688, 2856, 3024, 3192, 3360, 3528, 3696, 3864, 4032, 4200, 4368, 4536, 4704, 4872, 5040, 5208, 5376, 5544, 5712, 5880, 6048, 6216, 6384, 6552, 6720, 6888, 7056, 7224, 7392, 7560, 7728, 7896, 8064, 8232, 8400, 8568, 8736, 8904, 9072, 9240, 9408, 9576, 9744, 9912, 10080, 10248, 10416, 10584, 10752, 10920, 11088, 11256, 11424, 11592, 11760, 11928, 12096, 12264, 12432, 12600, 12768, 12936, 13104, 13272, 13440, 13608, 13776, 13944, 14112, 14280, 14448, 14616, 14784, 14952, 15120, 15288, 15456, 15624, 15792, 15960, 16128, 16296, 16464, 16632, 16800, 16968, 17136, 17304, 17472, 17640, 17808, 17976, 18144, 18312, 18480, 18648, 18816, 18984, 19152, 19320, 19488, 19656, 19824, 19992, 20160, 20328, 20496, 20664, 20832, 21000, 21168, 21336, 21504, 21672, 21840, 22008, 22176, 22344, 22512, 22680, 22848, 23016, 23184, 23352, 23520, 23688, 23856, 24024, 24192, 24360, 24528, 24696, 24864, 25032, 25200, 25368, 25536, 25704, 25872, 26040, 26208, 26376, 26544, 26712, 26880, 27048, 27216, 27384, 27552, 27720, 27888, 28056, 28224, 28392, 28560, 28728, 28896, 29064, 29232, 29400, 29568, 29736, 29904, 30072, 30240, 30408, 30576, 30744, 30912, 31080, 31248, 31416, 31584, 31752, 31920, 32088, 32256, 32424, 32592, 32760, 32928, 33096, 33264, 33432, 33600, 33768, 33936, 34104, 34272, 34440, 34608, 34776, 34944, 35112, 35280, 35448, 35616, 35784, 35952, 36120, 36288, 36456, 36624, 36792, 36960, 37128, 37296, 37464, 37632, 37800, 37968, 38136, 38304, 38472, 38640, 38808, 38976, 39144, 39312, 39480, 39648, 39816, 39984, 40152, 40320, 40488, 40656, 40824, 40992, 41160, 41328, 41496, 41664, 41832, 42000, 42168, 42336, 42504, 42672, 42840, 
0, 169, 338, 507, 676, 845, 1014, 1183, 1352, 1521, 1690, 1859, 2028, 2197, 2366, 2535, 2704, 2873, 3042, 3211, 3380, 3549, 3718, 3887, 4056, 4225, 4394, 4563, 4732, 4901, 5070, 5239, 5408, 5577, 5746, 5915, 6084, 6253, 6422, 6591, 6760, 6929, 7098, 7267, 7436, 7605, 7774, 7943, 8112, 8281, 8450, 8619, 8788, 8957, 9126, 9295, 9464, 9633, 9802, 9971, 10140, 10309, 10478, 10647, 10816, 10985, 11154, 11323, 11492, 11661, 11830, 11999, 12168, 12337, 12506, 12675, 12844, 13013, 13182, 13351, 13520, 13689, 13858, 14027, 14196, 14365, 14534, 14703, 14872, 15041, 15210, 15379, 15548, 15717, 15886, 16055, 16224, 16393, 16562, 16731, 16900, 17069, 17238, 17407, 17576, 17745, 17914, 18083, 18252, 18421, 18590, 18759, 18928, 19097, 19266, 19435, 19604, 19773, 19942, 20111, 20280, 20449, 20618, 20787, 20956, 21125, 21294, 21463, 21632, 21801, 21970, 22139, 22308, 22477, 22646, 22815, 22984, 23153, 23322, 23491, 23660, 23829, 23998, 24167, 24336, 24505, 24674, 24843, 25012, 25181, 25350, 25519, 25688, 25857, 26026, 26195, 26364, 26533, 26702, 26871, 27040, 27209, 27378, 27547, 27716, 27885, 28054, 28223, 28392, 28561, 28730, 28899, 29068, 29237, 29406, 29575, 29744, 29913, 30082, 30251, 30420, 30589, 30758, 30927, 31096, 31265, 31434, 31603, 31772, 31941, 32110, 32279, 32448, 32617, 32786, 32955, 33124, 33293, 33462, 33631, 33800, 33969, 34138, 34307, 34476, 34645, 34814, 34983, 35152, 35321, 35490, 35659, 35828, 35997, 36166, 36335, 36504, 36673, 36842, 37011, 37180, 37349, 37518, 37687, 37856, 38025, 38194, 38363, 38532, 38701, 38870, 39039, 39208, 39377, 39546, 39715, 39884, 40053, 40222, 40391, 40560, 40729, 40898, 41067, 41236, 41405, 41574, 41743, 41912, 42081, 42250, 42419, 42588, 42757, 42926, 43095, 
0, 170, 340, 510, 680, 850, 1020, 1190, 1360, 1530, 1700, 1870, 2040, 2210, 2380, 2550, 2720, 2890, 3060, 3230, 3400, 3570, 3740, 3910, 4080, 4250, 4420, 4590, 4760, 4930, 5100, 5270, 5440, 5610, 5780, 5950, 6120, 6290, 6460, 6630, 6800, 6970, 7140, 7310, 7480, 7650, 7820, 7990, 8160, 8330, 8500, 8670, 8840, 9010, 9180, 9350, 9520, 9690, 9860, 10030, 10200, 10370, 10540, 10710, 10880, 11050, 11220, 11390, 11560, 11730, 11900, 12070, 12240, 12410, 12580, 12750, 12920, 13090, 13260, 13430, 13600, 13770, 13940, 14110, 14280, 14450, 14620, 14790, 14960, 15130, 15300, 15470, 15640, 15810, 15980, 16150, 16320, 16490, 16660, 16830, 17000, 17170, 17340, 17510, 17680, 17850, 18020, 18190, 18360, 18530, 18700, 18870, 19040, 19210, 19380, 19550, 19720, 19890, 20060, 20230, 20400, 20570, 20740, 20910, 21080, 21250, 21420, 21590, 21760, 21930, 22100, 22270, 22440, 22610, 22780, 22950, 23120, 23290, 23460, 23630, 23800, 23970, 24140, 24310, 24480, 24650, 24820, 24990, 25160, 25330, 25500, 25670, 25840, 26010, 26180, 26350, 26520, 26690, 26860, 27030, 27200, 27370, 27540, 27710, 27880, 28050, 28220, 28390, 28560, 28730, 28900, 29070, 29240, 29410, 29580, 29750, 29920, 30090, 30260, 30430, 30600, 30770, 30940, 31110, 31280, 31450, 31620, 31790, 31960, 32130, 32300, 32470, 32640, 32810, 32980, 33150, 33320, 33490, 33660, 33830, 34000, 34170, 34340, 34510, 34680, 34850, 35020, 35190, 35360, 35530, 35700, 35870, 36040, 36210, 36380, 36550, 36720, 36890, 37060, 37230, 37400, 37570, 37740, 37910, 38080, 38250, 38420, 38590, 38760, 38930, 39100, 39270, 39440, 39610, 39780, 39950, 40120, 40290, 40460, 40630, 40800, 40970, 41140, 41310, 41480, 41650, 41820, 41990, 42160, 42330, 42500, 42670, 42840, 43010, 43180, 43350, 
0, 171, 342, 513, 684, 855, 1026, 1197, 1368, 1539, 1710, 1881, 2052, 2223, 2394, 2565, 2736, 2907, 3078, 3249, 3420, 3591, 3762, 3933, 4104, 4275, 4446, 4617, 4788, 4959, 5130, 5301, 5472, 5643, 5814, 5985, 6156, 6327, 6498, 6669, 6840, 7011, 7182, 7353, 7524, 7695, 7866, 8037, 8208, 8379, 8550, 8721, 8892, 9063, 9234, 9405, 9576, 9747, 9918, 10089, 10260, 10431, 10602, 10773, 10944, 11115, 11286, 11457, 11628, 11799, 11970, 12141, 12312, 12483, 12654, 12825, 12996, 13167, 13338, 13509, 13680, 13851, 14022, 14193, 14364, 14535, 14706, 14877, 15048, 15219, 15390, 15561, 15732, 15903, 16074, 16245, 16416, 16587, 16758, 16929, 17100, 17271, 17442, 17613, 17784, 17955, 18126, 18297, 18468, 18639, 18810, 18981, 19152, 19323, 19494, 19665, 19836, 20007, 20178, 20349, 20520, 20691, 20862, 21033, 21204, 21375, 21546, 21717, 21888, 22059, 22230, 22401, 22572, 22743, 22914, 23085, 23256, 23427, 23598, 23769, 23940, 24111, 24282, 24453, 24624, 24795, 24966, 25137, 25308, 25479, 25650, 25821, 25992, 26163, 26334, 26505, 26676, 26847, 27018, 27189, 27360, 27531, 27702, 27873, 28044, 28215, 28386, 28557, 28728, 28899, 29070, 29241, 29412, 29583, 29754, 29925, 30096, 30267, 30438, 30609, 30780, 30951, 31122, 31293, 31464, 31635, 31806, 31977, 32148, 32319, 32490, 32661, 32832, 33003, 33174, 33345, 33516, 33687, 33858, 34029, 34200, 34371, 34542, 34713, 34884, 35055, 35226, 35397, 35568, 35739, 35910, 36081, 36252, 36423, 36594, 36765, 36936, 37107, 37278, 37449, 37620, 37791, 37962, 38133, 38304, 38475, 38646, 38817, 38988, 39159, 39330, 39501, 39672, 39843, 40014, 40185, 40356, 40527, 40698, 40869, 41040, 41211, 41382, 41553, 41724, 41895, 42066, 42237, 42408, 42579, 42750, 42921, 43092, 43263, 43434, 43605, 
0, 172, 344, 516, 688, 860, 1032, 1204, 1376, 1548, 1720, 1892, 2064, 2236, 2408, 2580, 2752, 2924, 3096, 3268, 3440, 3612, 3784, 3956, 4128, 4300, 4472, 4644, 4816, 4988, 5160, 5332, 5504, 5676, 5848, 6020, 6192, 6364, 6536, 6708, 6880, 7052, 7224, 7396, 7568, 7740, 7912, 8084, 8256, 8428, 8600, 8772, 8944, 9116, 9288, 9460, 9632, 9804, 9976, 10148, 10320, 10492, 10664, 10836, 11008, 11180, 11352, 11524, 11696, 11868, 12040, 12212, 12384, 12556, 12728, 12900, 13072, 13244, 13416, 13588, 13760, 13932, 14104, 14276, 14448, 14620, 14792, 14964, 15136, 15308, 15480, 15652, 15824, 15996, 16168, 16340, 16512, 16684, 16856, 17028, 17200, 17372, 17544, 17716, 17888, 18060, 18232, 18404, 18576, 18748, 18920, 19092, 19264, 19436, 19608, 19780, 19952, 20124, 20296, 20468, 20640, 20812, 20984, 21156, 21328, 21500, 21672, 21844, 22016, 22188, 22360, 22532, 22704, 22876, 23048, 23220, 23392, 23564, 23736, 23908, 24080, 24252, 24424, 24596, 24768, 24940, 25112, 25284, 25456, 25628, 25800, 25972, 26144, 26316, 26488, 26660, 26832, 27004, 27176, 27348, 27520, 27692, 27864, 28036, 28208, 28380, 28552, 28724, 28896, 29068, 29240, 29412, 29584, 29756, 29928, 30100, 30272, 30444, 30616, 30788, 30960, 31132, 31304, 31476, 31648, 31820, 31992, 32164, 32336, 32508, 32680, 32852, 33024, 33196, 33368, 33540, 33712, 33884, 34056, 34228, 34400, 34572, 34744, 34916, 35088, 35260, 35432, 35604, 35776, 35948, 36120, 36292, 36464, 36636, 36808, 36980, 37152, 37324, 37496, 37668, 37840, 38012, 38184, 38356, 38528, 38700, 38872, 39044, 39216, 39388, 39560, 39732, 39904, 40076, 40248, 40420, 40592, 40764, 40936, 41108, 41280, 41452, 41624, 41796, 41968, 42140, 42312, 42484, 42656, 42828, 43000, 43172, 43344, 43516, 43688, 43860, 
0, 173, 346, 519, 692, 865, 1038, 1211, 1384, 1557, 1730, 1903, 2076, 2249, 2422, 2595, 2768, 2941, 3114, 3287, 3460, 3633, 3806, 3979, 4152, 4325, 4498, 4671, 4844, 5017, 5190, 5363, 5536, 5709, 5882, 6055, 6228, 6401, 6574, 6747, 6920, 7093, 7266, 7439, 7612, 7785, 7958, 8131, 8304, 8477, 8650, 8823, 8996, 9169, 9342, 9515, 9688, 9861, 10034, 10207, 10380, 10553, 10726, 10899, 11072, 11245, 11418, 11591, 11764, 11937, 12110, 12283, 12456, 12629, 12802, 12975, 13148, 13321, 13494, 13667, 13840, 14013, 14186, 14359, 14532, 14705, 14878, 15051, 15224, 15397, 15570, 15743, 15916, 16089, 16262, 16435, 16608, 16781, 16954, 17127, 17300, 17473, 17646, 17819, 17992, 18165, 18338, 18511, 18684, 18857, 19030, 19203, 19376, 19549, 19722, 19895, 20068, 20241, 20414, 20587, 20760, 20933, 21106, 21279, 21452, 21625, 21798, 21971, 22144, 22317, 22490, 22663, 22836, 23009, 23182, 23355, 23528, 23701, 23874, 24047, 24220, 24393, 24566, 24739, 24912, 25085, 25258, 25431, 25604, 25777, 25950, 26123, 26296, 26469, 26642, 26815, 26988, 27161, 27334, 27507, 27680, 27853, 28026, 28199, 28372, 28545, 28718, 28891, 29064, 29237, 29410, 29583, 29756, 29929, 30102, 30275, 30448, 30621, 30794, 30967, 31140, 31313, 31486, 31659, 31832, 32005, 32178, 32351, 32524, 32697, 32870, 33043, 33216, 33389, 33562, 33735, 33908, 34081, 34254, 34427, 34600, 34773, 34946, 35119, 35292, 35465, 35638, 35811, 35984, 36157, 36330, 36503, 36676, 36849, 37022, 37195, 37368, 37541, 37714, 37887, 38060, 38233, 38406, 38579, 38752, 38925, 39098, 39271, 39444, 39617, 39790, 39963, 40136, 40309, 40482, 40655, 40828, 41001, 41174, 41347, 41520, 41693, 41866, 42039, 42212, 42385, 42558, 42731, 42904, 43077, 43250, 43423, 43596, 43769, 43942, 44115, 
0, 174, 348, 522, 696, 870, 1044, 1218, 1392, 1566, 1740, 1914, 2088, 2262, 2436, 2610, 2784, 2958, 3132, 3306, 3480, 3654, 3828, 4002, 4176, 4350, 4524, 4698, 4872, 5046, 5220, 5394, 5568, 5742, 5916, 6090, 6264, 6438, 6612, 6786, 6960, 7134, 7308, 7482, 7656, 7830, 8004, 8178, 8352, 8526, 8700, 8874, 9048, 9222, 9396, 9570, 9744, 9918, 10092, 10266, 10440, 10614, 10788, 10962, 11136, 11310, 11484, 11658, 11832, 12006, 12180, 12354, 12528, 12702, 12876, 13050, 13224, 13398, 13572, 13746, 13920, 14094, 14268, 14442, 14616, 14790, 14964, 15138, 15312, 15486, 15660, 15834, 16008, 16182, 16356, 16530, 16704, 16878, 17052, 17226, 17400, 17574, 17748, 17922, 18096, 18270, 18444, 18618, 18792, 18966, 19140, 19314, 19488, 19662, 19836, 20010, 20184, 20358, 20532, 20706, 20880, 21054, 21228, 21402, 21576, 21750, 21924, 22098, 22272, 22446, 22620, 22794, 22968, 23142, 23316, 23490, 23664, 23838, 24012, 24186, 24360, 24534, 24708, 24882, 25056, 25230, 25404, 25578, 25752, 25926, 26100, 26274, 26448, 26622, 26796, 26970, 27144, 27318, 27492, 27666, 27840, 28014, 28188, 28362, 28536, 28710, 28884, 29058, 29232, 29406, 29580, 29754, 29928, 30102, 30276, 30450, 30624, 30798, 30972, 31146, 31320, 31494, 31668, 31842, 32016, 32190, 32364, 32538, 32712, 32886, 33060, 33234, 33408, 33582, 33756, 33930, 34104, 34278, 34452, 34626, 34800, 34974, 35148, 35322, 35496, 35670, 35844, 36018, 36192, 36366, 36540, 36714, 36888, 37062, 37236, 37410, 37584, 37758, 37932, 38106, 38280, 38454, 38628, 38802, 38976, 39150, 39324, 39498, 39672, 39846, 40020, 40194, 40368, 40542, 40716, 40890, 41064, 41238, 41412, 41586, 41760, 41934, 42108, 42282, 42456, 42630, 42804, 42978, 43152, 43326, 43500, 43674, 43848, 44022, 44196, 44370, 
0, 175, 350, 525, 700, 875, 1050, 1225, 1400, 1575, 1750, 1925, 2100, 2275, 2450, 2625, 2800, 2975, 3150, 3325, 3500, 3675, 3850, 4025, 4200, 4375, 4550, 4725, 4900, 5075, 5250, 5425, 5600, 5775, 5950, 6125, 6300, 6475, 6650, 6825, 7000, 7175, 7350, 7525, 7700, 7875, 8050, 8225, 8400, 8575, 8750, 8925, 9100, 9275, 9450, 9625, 9800, 9975, 10150, 10325, 10500, 10675, 10850, 11025, 11200, 11375, 11550, 11725, 11900, 12075, 12250, 12425, 12600, 12775, 12950, 13125, 13300, 13475, 13650, 13825, 14000, 14175, 14350, 14525, 14700, 14875, 15050, 15225, 15400, 15575, 15750, 15925, 16100, 16275, 16450, 16625, 16800, 16975, 17150, 17325, 17500, 17675, 17850, 18025, 18200, 18375, 18550, 18725, 18900, 19075, 19250, 19425, 19600, 19775, 19950, 20125, 20300, 20475, 20650, 20825, 21000, 21175, 21350, 21525, 21700, 21875, 22050, 22225, 22400, 22575, 22750, 22925, 23100, 23275, 23450, 23625, 23800, 23975, 24150, 24325, 24500, 24675, 24850, 25025, 25200, 25375, 25550, 25725, 25900, 26075, 26250, 26425, 26600, 26775, 26950, 27125, 27300, 27475, 27650, 27825, 28000, 28175, 28350, 28525, 28700, 28875, 29050, 29225, 29400, 29575, 29750, 29925, 30100, 30275, 30450, 30625, 30800, 30975, 31150, 31325, 31500, 31675, 31850, 32025, 32200, 32375, 32550, 32725, 32900, 33075, 33250, 33425, 33600, 33775, 33950, 34125, 34300, 34475, 34650, 34825, 35000, 35175, 35350, 35525, 35700, 35875, 36050, 36225, 36400, 36575, 36750, 36925, 37100, 37275, 37450, 37625, 37800, 37975, 38150, 38325, 38500, 38675, 38850, 39025, 39200, 39375, 39550, 39725, 39900, 40075, 40250, 40425, 40600, 40775, 40950, 41125, 41300, 41475, 41650, 41825, 42000, 42175, 42350, 42525, 42700, 42875, 43050, 43225, 43400, 43575, 43750, 43925, 44100, 44275, 44450, 44625, 
0, 176, 352, 528, 704, 880, 1056, 1232, 1408, 1584, 1760, 1936, 2112, 2288, 2464, 2640, 2816, 2992, 3168, 3344, 3520, 3696, 3872, 4048, 4224, 4400, 4576, 4752, 4928, 5104, 5280, 5456, 5632, 5808, 5984, 6160, 6336, 6512, 6688, 6864, 7040, 7216, 7392, 7568, 7744, 7920, 8096, 8272, 8448, 8624, 8800, 8976, 9152, 9328, 9504, 9680, 9856, 10032, 10208, 10384, 10560, 10736, 10912, 11088, 11264, 11440, 11616, 11792, 11968, 12144, 12320, 12496, 12672, 12848, 13024, 13200, 13376, 13552, 13728, 13904, 14080, 14256, 14432, 14608, 14784, 14960, 15136, 15312, 15488, 15664, 15840, 16016, 16192, 16368, 16544, 16720, 16896, 17072, 17248, 17424, 17600, 17776, 17952, 18128, 18304, 18480, 18656, 18832, 19008, 19184, 19360, 19536, 19712, 19888, 20064, 20240, 20416, 20592, 20768, 20944, 21120, 21296, 21472, 21648, 21824, 22000, 22176, 22352, 22528, 22704, 22880, 23056, 23232, 23408, 23584, 23760, 23936, 24112, 24288, 24464, 24640, 24816, 24992, 25168, 25344, 25520, 25696, 25872, 26048, 26224, 26400, 26576, 26752, 26928, 27104, 27280, 27456, 27632, 27808, 27984, 28160, 28336, 28512, 28688, 28864, 29040, 29216, 29392, 29568, 29744, 29920, 30096, 30272, 30448, 30624, 30800, 30976, 31152, 31328, 31504, 31680, 31856, 32032, 32208, 32384, 32560, 32736, 32912, 33088, 33264, 33440, 33616, 33792, 33968, 34144, 34320, 34496, 34672, 34848, 35024, 35200, 35376, 35552, 35728, 35904, 36080, 36256, 36432, 36608, 36784, 36960, 37136, 37312, 37488, 37664, 37840, 38016, 38192, 38368, 38544, 38720, 38896, 39072, 39248, 39424, 39600, 39776, 39952, 40128, 40304, 40480, 40656, 40832, 41008, 41184, 41360, 41536, 41712, 41888, 42064, 42240, 42416, 42592, 42768, 42944, 43120, 43296, 43472, 43648, 43824, 44000, 44176, 44352, 44528, 44704, 44880, 
0, 177, 354, 531, 708, 885, 1062, 1239, 1416, 1593, 1770, 1947, 2124, 2301, 2478, 2655, 2832, 3009, 3186, 3363, 3540, 3717, 3894, 4071, 4248, 4425, 4602, 4779, 4956, 5133, 5310, 5487, 5664, 5841, 6018, 6195, 6372, 6549, 6726, 6903, 7080, 7257, 7434, 7611, 7788, 7965, 8142, 8319, 8496, 8673, 8850, 9027, 9204, 9381, 9558, 9735, 9912, 10089, 10266, 10443, 10620, 10797, 10974, 11151, 11328, 11505, 11682, 11859, 12036, 12213, 12390, 12567, 12744, 12921, 13098, 13275, 13452, 13629, 13806, 13983, 14160, 14337, 14514, 14691, 14868, 15045, 15222, 15399, 15576, 15753, 15930, 16107, 16284, 16461, 16638, 16815, 16992, 17169, 17346, 17523, 17700, 17877, 18054, 18231, 18408, 18585, 18762, 18939, 19116, 19293, 19470, 19647, 19824, 20001, 20178, 20355, 20532, 20709, 20886, 21063, 21240, 21417, 21594, 21771, 21948, 22125, 22302, 22479, 22656, 22833, 23010, 23187, 23364, 23541, 23718, 23895, 24072, 24249, 24426, 24603, 24780, 24957, 25134, 25311, 25488, 25665, 25842, 26019, 26196, 26373, 26550, 26727, 26904, 27081, 27258, 27435, 27612, 27789, 27966, 28143, 28320, 28497, 28674, 28851, 29028, 29205, 29382, 29559, 29736, 29913, 30090, 30267, 30444, 30621, 30798, 30975, 31152, 31329, 31506, 31683, 31860, 32037, 32214, 32391, 32568, 32745, 32922, 33099, 33276, 33453, 33630, 33807, 33984, 34161, 34338, 34515, 34692, 34869, 35046, 35223, 35400, 35577, 35754, 35931, 36108, 36285, 36462, 36639, 36816, 36993, 37170, 37347, 37524, 37701, 37878, 38055, 38232, 38409, 38586, 38763, 38940, 39117, 39294, 39471, 39648, 39825, 40002, 40179, 40356, 40533, 40710, 40887, 41064, 41241, 41418, 41595, 41772, 41949, 42126, 42303, 42480, 42657, 42834, 43011, 43188, 43365, 43542, 43719, 43896, 44073, 44250, 44427, 44604, 44781, 44958, 45135, 
0, 178, 356, 534, 712, 890, 1068, 1246, 1424, 1602, 1780, 1958, 2136, 2314, 2492, 2670, 2848, 3026, 3204, 3382, 3560, 3738, 3916, 4094, 4272, 4450, 4628, 4806, 4984, 5162, 5340, 5518, 5696, 5874, 6052, 6230, 6408, 6586, 6764, 6942, 7120, 7298, 7476, 7654, 7832, 8010, 8188, 8366, 8544, 8722, 8900, 9078, 9256, 9434, 9612, 9790, 9968, 10146, 10324, 10502, 10680, 10858, 11036, 11214, 11392, 11570, 11748, 11926, 12104, 12282, 12460, 12638, 12816, 12994, 13172, 13350, 13528, 13706, 13884, 14062, 14240, 14418, 14596, 14774, 14952, 15130, 15308, 15486, 15664, 15842, 16020, 16198, 16376, 16554, 16732, 16910, 17088, 17266, 17444, 17622, 17800, 17978, 18156, 18334, 18512, 18690, 18868, 19046, 19224, 19402, 19580, 19758, 19936, 20114, 20292, 20470, 20648, 20826, 21004, 21182, 21360, 21538, 21716, 21894, 22072, 22250, 22428, 22606, 22784, 22962, 23140, 23318, 23496, 23674, 23852, 24030, 24208, 24386, 24564, 24742, 24920, 25098, 25276, 25454, 25632, 25810, 25988, 26166, 26344, 26522, 26700, 26878, 27056, 27234, 27412, 27590, 27768, 27946, 28124, 28302, 28480, 28658, 28836, 29014, 29192, 29370, 29548, 29726, 29904, 30082, 30260, 30438, 30616, 30794, 30972, 31150, 31328, 31506, 31684, 31862, 32040, 32218, 32396, 32574, 32752, 32930, 33108, 33286, 33464, 33642, 33820, 33998, 34176, 34354, 34532, 34710, 34888, 35066, 35244, 35422, 35600, 35778, 35956, 36134, 36312, 36490, 36668, 36846, 37024, 37202, 37380, 37558, 37736, 37914, 38092, 38270, 38448, 38626, 38804, 38982, 39160, 39338, 39516, 39694, 39872, 40050, 40228, 40406, 40584, 40762, 40940, 41118, 41296, 41474, 41652, 41830, 42008, 42186, 42364, 42542, 42720, 42898, 43076, 43254, 43432, 43610, 43788, 43966, 44144, 44322, 44500, 44678, 44856, 45034, 45212, 45390, 
0, 179, 358, 537, 716, 895, 1074, 1253, 1432, 1611, 1790, 1969, 2148, 2327, 2506, 2685, 2864, 3043, 3222, 3401, 3580, 3759, 3938, 4117, 4296, 4475, 4654, 4833, 5012, 5191, 5370, 5549, 5728, 5907, 6086, 6265, 6444, 6623, 6802, 6981, 7160, 7339, 7518, 7697, 7876, 8055, 8234, 8413, 8592, 8771, 8950, 9129, 9308, 9487, 9666, 9845, 10024, 10203, 10382, 10561, 10740, 10919, 11098, 11277, 11456, 11635, 11814, 11993, 12172, 12351, 12530, 12709, 12888, 13067, 13246, 13425, 13604, 13783, 13962, 14141, 14320, 14499, 14678, 14857, 15036, 15215, 15394, 15573, 15752, 15931, 16110, 16289, 16468, 16647, 16826, 17005, 17184, 17363, 17542, 17721, 17900, 18079, 18258, 18437, 18616, 18795, 18974, 19153, 19332, 19511, 19690, 19869, 20048, 20227, 20406, 20585, 20764, 20943, 21122, 21301, 21480, 21659, 21838, 22017, 22196, 22375, 22554, 22733, 22912, 23091, 23270, 23449, 23628, 23807, 23986, 24165, 24344, 24523, 24702, 24881, 25060, 25239, 25418, 25597, 25776, 25955, 26134, 26313, 26492, 26671, 26850, 27029, 27208, 27387, 27566, 27745, 27924, 28103, 28282, 28461, 28640, 28819, 28998, 29177, 29356, 29535, 29714, 29893, 30072, 30251, 30430, 30609, 30788, 30967, 31146, 31325, 31504, 31683, 31862, 32041, 32220, 32399, 32578, 32757, 32936, 33115, 33294, 33473, 33652, 33831, 34010, 34189, 34368, 34547, 34726, 34905, 35084, 35263, 35442, 35621, 35800, 35979, 36158, 36337, 36516, 36695, 36874, 37053, 37232, 37411, 37590, 37769, 37948, 38127, 38306, 38485, 38664, 38843, 39022, 39201, 39380, 39559, 39738, 39917, 40096, 40275, 40454, 40633, 40812, 40991, 41170, 41349, 41528, 41707, 41886, 42065, 42244, 42423, 42602, 42781, 42960, 43139, 43318, 43497, 43676, 43855, 44034, 44213, 44392, 44571, 44750, 44929, 45108, 45287, 45466, 45645, 
0, 180, 360, 540, 720, 900, 1080, 1260, 1440, 1620, 1800, 1980, 2160, 2340, 2520, 2700, 2880, 3060, 3240, 3420, 3600, 3780, 3960, 4140, 4320, 4500, 4680, 4860, 5040, 5220, 5400, 5580, 5760, 5940, 6120, 6300, 6480, 6660, 6840, 7020, 7200, 7380, 7560, 7740, 7920, 8100, 8280, 8460, 8640, 8820, 9000, 9180, 9360, 9540, 9720, 9900, 10080, 10260, 10440, 10620, 10800, 10980, 11160, 11340, 11520, 11700, 11880, 12060, 12240, 12420, 12600, 12780, 12960, 13140, 13320, 13500, 13680, 13860, 14040, 14220, 14400, 14580, 14760, 14940, 15120, 15300, 15480, 15660, 15840, 16020, 16200, 16380, 16560, 16740, 16920, 17100, 17280, 17460, 17640, 17820, 18000, 18180, 18360, 18540, 18720, 18900, 19080, 19260, 19440, 19620, 19800, 19980, 20160, 20340, 20520, 20700, 20880, 21060, 21240, 21420, 21600, 21780, 21960, 22140, 22320, 22500, 22680, 22860, 23040, 23220, 23400, 23580, 23760, 23940, 24120, 24300, 24480, 24660, 24840, 25020, 25200, 25380, 25560, 25740, 25920, 26100, 26280, 26460, 26640, 26820, 27000, 27180, 27360, 27540, 27720, 27900, 28080, 28260, 28440, 28620, 28800, 28980, 29160, 29340, 29520, 29700, 29880, 30060, 30240, 30420, 30600, 30780, 30960, 31140, 31320, 31500, 31680, 31860, 32040, 32220, 32400, 32580, 32760, 32940, 33120, 33300, 33480, 33660, 33840, 34020, 34200, 34380, 34560, 34740, 34920, 35100, 35280, 35460, 35640, 35820, 36000, 36180, 36360, 36540, 36720, 36900, 37080, 37260, 37440, 37620, 37800, 37980, 38160, 38340, 38520, 38700, 38880, 39060, 39240, 39420, 39600, 39780, 39960, 40140, 40320, 40500, 40680, 40860, 41040, 41220, 41400, 41580, 41760, 41940, 42120, 42300, 42480, 42660, 42840, 43020, 43200, 43380, 43560, 43740, 43920, 44100, 44280, 44460, 44640, 44820, 45000, 45180, 45360, 45540, 45720, 45900, 
0, 181, 362, 543, 724, 905, 1086, 1267, 1448, 1629, 1810, 1991, 2172, 2353, 2534, 2715, 2896, 3077, 3258, 3439, 3620, 3801, 3982, 4163, 4344, 4525, 4706, 4887, 5068, 5249, 5430, 5611, 5792, 5973, 6154, 6335, 6516, 6697, 6878, 7059, 7240, 7421, 7602, 7783, 7964, 8145, 8326, 8507, 8688, 8869, 9050, 9231, 9412, 9593, 9774, 9955, 10136, 10317, 10498, 10679, 10860, 11041, 11222, 11403, 11584, 11765, 11946, 12127, 12308, 12489, 12670, 12851, 13032, 13213, 13394, 13575, 13756, 13937, 14118, 14299, 14480, 14661, 14842, 15023, 15204, 15385, 15566, 15747, 15928, 16109, 16290, 16471, 16652, 16833, 17014, 17195, 17376, 17557, 17738, 17919, 18100, 18281, 18462, 18643, 18824, 19005, 19186, 19367, 19548, 19729, 19910, 20091, 20272, 20453, 20634, 20815, 20996, 21177, 21358, 21539, 21720, 21901, 22082, 22263, 22444, 22625, 22806, 22987, 23168, 23349, 23530, 23711, 23892, 24073, 24254, 24435, 24616, 24797, 24978, 25159, 25340, 25521, 25702, 25883, 26064, 26245, 26426, 26607, 26788, 26969, 27150, 27331, 27512, 27693, 27874, 28055, 28236, 28417, 28598, 28779, 28960, 29141, 29322, 29503, 29684, 29865, 30046, 30227, 30408, 30589, 30770, 30951, 31132, 31313, 31494, 31675, 31856, 32037, 32218, 32399, 32580, 32761, 32942, 33123, 33304, 33485, 33666, 33847, 34028, 34209, 34390, 34571, 34752, 34933, 35114, 35295, 35476, 35657, 35838, 36019, 36200, 36381, 36562, 36743, 36924, 37105, 37286, 37467, 37648, 37829, 38010, 38191, 38372, 38553, 38734, 38915, 39096, 39277, 39458, 39639, 39820, 40001, 40182, 40363, 40544, 40725, 40906, 41087, 41268, 41449, 41630, 41811, 41992, 42173, 42354, 42535, 42716, 42897, 43078, 43259, 43440, 43621, 43802, 43983, 44164, 44345, 44526, 44707, 44888, 45069, 45250, 45431, 45612, 45793, 45974, 46155, 
0, 182, 364, 546, 728, 910, 1092, 1274, 1456, 1638, 1820, 2002, 2184, 2366, 2548, 2730, 2912, 3094, 3276, 3458, 3640, 3822, 4004, 4186, 4368, 4550, 4732, 4914, 5096, 5278, 5460, 5642, 5824, 6006, 6188, 6370, 6552, 6734, 6916, 7098, 7280, 7462, 7644, 7826, 8008, 8190, 8372, 8554, 8736, 8918, 9100, 9282, 9464, 9646, 9828, 10010, 10192, 10374, 10556, 10738, 10920, 11102, 11284, 11466, 11648, 11830, 12012, 12194, 12376, 12558, 12740, 12922, 13104, 13286, 13468, 13650, 13832, 14014, 14196, 14378, 14560, 14742, 14924, 15106, 15288, 15470, 15652, 15834, 16016, 16198, 16380, 16562, 16744, 16926, 17108, 17290, 17472, 17654, 17836, 18018, 18200, 18382, 18564, 18746, 18928, 19110, 19292, 19474, 19656, 19838, 20020, 20202, 20384, 20566, 20748, 20930, 21112, 21294, 21476, 21658, 21840, 22022, 22204, 22386, 22568, 22750, 22932, 23114, 23296, 23478, 23660, 23842, 24024, 24206, 24388, 24570, 24752, 24934, 25116, 25298, 25480, 25662, 25844, 26026, 26208, 26390, 26572, 26754, 26936, 27118, 27300, 27482, 27664, 27846, 28028, 28210, 28392, 28574, 28756, 28938, 29120, 29302, 29484, 29666, 29848, 30030, 30212, 30394, 30576, 30758, 30940, 31122, 31304, 31486, 31668, 31850, 32032, 32214, 32396, 32578, 32760, 32942, 33124, 33306, 33488, 33670, 33852, 34034, 34216, 34398, 34580, 34762, 34944, 35126, 35308, 35490, 35672, 35854, 36036, 36218, 36400, 36582, 36764, 36946, 37128, 37310, 37492, 37674, 37856, 38038, 38220, 38402, 38584, 38766, 38948, 39130, 39312, 39494, 39676, 39858, 40040, 40222, 40404, 40586, 40768, 40950, 41132, 41314, 41496, 41678, 41860, 42042, 42224, 42406, 42588, 42770, 42952, 43134, 43316, 43498, 43680, 43862, 44044, 44226, 44408, 44590, 44772, 44954, 45136, 45318, 45500, 45682, 45864, 46046, 46228, 46410, 
0, 183, 366, 549, 732, 915, 1098, 1281, 1464, 1647, 1830, 2013, 2196, 2379, 2562, 2745, 2928, 3111, 3294, 3477, 3660, 3843, 4026, 4209, 4392, 4575, 4758, 4941, 5124, 5307, 5490, 5673, 5856, 6039, 6222, 6405, 6588, 6771, 6954, 7137, 7320, 7503, 7686, 7869, 8052, 8235, 8418, 8601, 8784, 8967, 9150, 9333, 9516, 9699, 9882, 10065, 10248, 10431, 10614, 10797, 10980, 11163, 11346, 11529, 11712, 11895, 12078, 12261, 12444, 12627, 12810, 12993, 13176, 13359, 13542, 13725, 13908, 14091, 14274, 14457, 14640, 14823, 15006, 15189, 15372, 15555, 15738, 15921, 16104, 16287, 16470, 16653, 16836, 17019, 17202, 17385, 17568, 17751, 17934, 18117, 18300, 18483, 18666, 18849, 19032, 19215, 19398, 19581, 19764, 19947, 20130, 20313, 20496, 20679, 20862, 21045, 21228, 21411, 21594, 21777, 21960, 22143, 22326, 22509, 22692, 22875, 23058, 23241, 23424, 23607, 23790, 23973, 24156, 24339, 24522, 24705, 24888, 25071, 25254, 25437, 25620, 25803, 25986, 26169, 26352, 26535, 26718, 26901, 27084, 27267, 27450, 27633, 27816, 27999, 28182, 28365, 28548, 28731, 28914, 29097, 29280, 29463, 29646, 29829, 30012, 30195, 30378, 30561, 30744, 30927, 31110, 31293, 31476, 31659, 31842, 32025, 32208, 32391, 32574, 32757, 32940, 33123, 33306, 33489, 33672, 33855, 34038, 34221, 34404, 34587, 34770, 34953, 35136, 35319, 35502, 35685, 35868, 36051, 36234, 36417, 36600, 36783, 36966, 37149, 37332, 37515, 37698, 37881, 38064, 38247, 38430, 38613, 38796, 38979, 39162, 39345, 39528, 39711, 39894, 40077, 40260, 40443, 40626, 40809, 40992, 41175, 41358, 41541, 41724, 41907, 42090, 42273, 42456, 42639, 42822, 43005, 43188, 43371, 43554, 43737, 43920, 44103, 44286, 44469, 44652, 44835, 45018, 45201, 45384, 45567, 45750, 45933, 46116, 46299, 46482, 46665, 
0, 184, 368, 552, 736, 920, 1104, 1288, 1472, 1656, 1840, 2024, 2208, 2392, 2576, 2760, 2944, 3128, 3312, 3496, 3680, 3864, 4048, 4232, 4416, 4600, 4784, 4968, 5152, 5336, 5520, 5704, 5888, 6072, 6256, 6440, 6624, 6808, 6992, 7176, 7360, 7544, 7728, 7912, 8096, 8280, 8464, 8648, 8832, 9016, 9200, 9384, 9568, 9752, 9936, 10120, 10304, 10488, 10672, 10856, 11040, 11224, 11408, 11592, 11776, 11960, 12144, 12328, 12512, 12696, 12880, 13064, 13248, 13432, 13616, 13800, 13984, 14168, 14352, 14536, 14720, 14904, 15088, 15272, 15456, 15640, 15824, 16008, 16192, 16376, 16560, 16744, 16928, 17112, 17296, 17480, 17664, 17848, 18032, 18216, 18400, 18584, 18768, 18952, 19136, 19320, 19504, 19688, 19872, 20056, 20240, 20424, 20608, 20792, 20976, 21160, 21344, 21528, 21712, 21896, 22080, 22264, 22448, 22632, 22816, 23000, 23184, 23368, 23552, 23736, 23920, 24104, 24288, 24472, 24656, 24840, 25024, 25208, 25392, 25576, 25760, 25944, 26128, 26312, 26496, 26680, 26864, 27048, 27232, 27416, 27600, 27784, 27968, 28152, 28336, 28520, 28704, 28888, 29072, 29256, 29440, 29624, 29808, 29992, 30176, 30360, 30544, 30728, 30912, 31096, 31280, 31464, 31648, 31832, 32016, 32200, 32384, 32568, 32752, 32936, 33120, 33304, 33488, 33672, 33856, 34040, 34224, 34408, 34592, 34776, 34960, 35144, 35328, 35512, 35696, 35880, 36064, 36248, 36432, 36616, 36800, 36984, 37168, 37352, 37536, 37720, 37904, 38088, 38272, 38456, 38640, 38824, 39008, 39192, 39376, 39560, 39744, 39928, 40112, 40296, 40480, 40664, 40848, 41032, 41216, 41400, 41584, 41768, 41952, 42136, 42320, 42504, 42688, 42872, 43056, 43240, 43424, 43608, 43792, 43976, 44160, 44344, 44528, 44712, 44896, 45080, 45264, 45448, 45632, 45816, 46000, 46184, 46368, 46552, 46736, 46920, 
0, 185, 370, 555, 740, 925, 1110, 1295, 1480, 1665, 1850, 2035, 2220, 2405, 2590, 2775, 2960, 3145, 3330, 3515, 3700, 3885, 4070, 4255, 4440, 4625, 4810, 4995, 5180, 5365, 5550, 5735, 5920, 6105, 6290, 6475, 6660, 6845, 7030, 7215, 7400, 7585, 7770, 7955, 8140, 8325, 8510, 8695, 8880, 9065, 9250, 9435, 9620, 9805, 9990, 10175, 10360, 10545, 10730, 10915, 11100, 11285, 11470, 11655, 11840, 12025, 12210, 12395, 12580, 12765, 12950, 13135, 13320, 13505, 13690, 13875, 14060, 14245, 14430, 14615, 14800, 14985, 15170, 15355, 15540, 15725, 15910, 16095, 16280, 16465, 16650, 16835, 17020, 17205, 17390, 17575, 17760, 17945, 18130, 18315, 18500, 18685, 18870, 19055, 19240, 19425, 19610, 19795, 19980, 20165, 20350, 20535, 20720, 20905, 21090, 21275, 21460, 21645, 21830, 22015, 22200, 22385, 22570, 22755, 22940, 23125, 23310, 23495, 23680, 23865, 24050, 24235, 24420, 24605, 24790, 24975, 25160, 25345, 25530, 25715, 25900, 26085, 26270, 26455, 26640, 26825, 27010, 27195, 27380, 27565, 27750, 27935, 28120, 28305, 28490, 28675, 28860, 29045, 29230, 29415, 29600, 29785, 29970, 30155, 30340, 30525, 30710, 30895, 31080, 31265, 31450, 31635, 31820, 32005, 32190, 32375, 32560, 32745, 32930, 33115, 33300, 33485, 33670, 33855, 34040, 34225, 34410, 34595, 34780, 34965, 35150, 35335, 35520, 35705, 35890, 36075, 36260, 36445, 36630, 36815, 37000, 37185, 37370, 37555, 37740, 37925, 38110, 38295, 38480, 38665, 38850, 39035, 39220, 39405, 39590, 39775, 39960, 40145, 40330, 40515, 40700, 40885, 41070, 41255, 41440, 41625, 41810, 41995, 42180, 42365, 42550, 42735, 42920, 43105, 43290, 43475, 43660, 43845, 44030, 44215, 44400, 44585, 44770, 44955, 45140, 45325, 45510, 45695, 45880, 46065, 46250, 46435, 46620, 46805, 46990, 47175, 
0, 186, 372, 558, 744, 930, 1116, 1302, 1488, 1674, 1860, 2046, 2232, 2418, 2604, 2790, 2976, 3162, 3348, 3534, 3720, 3906, 4092, 4278, 4464, 4650, 4836, 5022, 5208, 5394, 5580, 5766, 5952, 6138, 6324, 6510, 6696, 6882, 7068, 7254, 7440, 7626, 7812, 7998, 8184, 8370, 8556, 8742, 8928, 9114, 9300, 9486, 9672, 9858, 10044, 10230, 10416, 10602, 10788, 10974, 11160, 11346, 11532, 11718, 11904, 12090, 12276, 12462, 12648, 12834, 13020, 13206, 13392, 13578, 13764, 13950, 14136, 14322, 14508, 14694, 14880, 15066, 15252, 15438, 15624, 15810, 15996, 16182, 16368, 16554, 16740, 16926, 17112, 17298, 17484, 17670, 17856, 18042, 18228, 18414, 18600, 18786, 18972, 19158, 19344, 19530, 19716, 19902, 20088, 20274, 20460, 20646, 20832, 21018, 21204, 21390, 21576, 21762, 21948, 22134, 22320, 22506, 22692, 22878, 23064, 23250, 23436, 23622, 23808, 23994, 24180, 24366, 24552, 24738, 24924, 25110, 25296, 25482, 25668, 25854, 26040, 26226, 26412, 26598, 26784, 26970, 27156, 27342, 27528, 27714, 27900, 28086, 28272, 28458, 28644, 28830, 29016, 29202, 29388, 29574, 29760, 29946, 30132, 30318, 30504, 30690, 30876, 31062, 31248, 31434, 31620, 31806, 31992, 32178, 32364, 32550, 32736, 32922, 33108, 33294, 33480, 33666, 33852, 34038, 34224, 34410, 34596, 34782, 34968, 35154, 35340, 35526, 35712, 35898, 36084, 36270, 36456, 36642, 36828, 37014, 37200, 37386, 37572, 37758, 37944, 38130, 38316, 38502, 38688, 38874, 39060, 39246, 39432, 39618, 39804, 39990, 40176, 40362, 40548, 40734, 40920, 41106, 41292, 41478, 41664, 41850, 42036, 42222, 42408, 42594, 42780, 42966, 43152, 43338, 43524, 43710, 43896, 44082, 44268, 44454, 44640, 44826, 45012, 45198, 45384, 45570, 45756, 45942, 46128, 46314, 46500, 46686, 46872, 47058, 47244, 47430, 
0, 187, 374, 561, 748, 935, 1122, 1309, 1496, 1683, 1870, 2057, 2244, 2431, 2618, 2805, 2992, 3179, 3366, 3553, 3740, 3927, 4114, 4301, 4488, 4675, 4862, 5049, 5236, 5423, 5610, 5797, 5984, 6171, 6358, 6545, 6732, 6919, 7106, 7293, 7480, 7667, 7854, 8041, 8228, 8415, 8602, 8789, 8976, 9163, 9350, 9537, 9724, 9911, 10098, 10285, 10472, 10659, 10846, 11033, 11220, 11407, 11594, 11781, 11968, 12155, 12342, 12529, 12716, 12903, 13090, 13277, 13464, 13651, 13838, 14025, 14212, 14399, 14586, 14773, 14960, 15147, 15334, 15521, 15708, 15895, 16082, 16269, 16456, 16643, 16830, 17017, 17204, 17391, 17578, 17765, 17952, 18139, 18326, 18513, 18700, 18887, 19074, 19261, 19448, 19635, 19822, 20009, 20196, 20383, 20570, 20757, 20944, 21131, 21318, 21505, 21692, 21879, 22066, 22253, 22440, 22627, 22814, 23001, 23188, 23375, 23562, 23749, 23936, 24123, 24310, 24497, 24684, 24871, 25058, 25245, 25432, 25619, 25806, 25993, 26180, 26367, 26554, 26741, 26928, 27115, 27302, 27489, 27676, 27863, 28050, 28237, 28424, 28611, 28798, 28985, 29172, 29359, 29546, 29733, 29920, 30107, 30294, 30481, 30668, 30855, 31042, 31229, 31416, 31603, 31790, 31977, 32164, 32351, 32538, 32725, 32912, 33099, 33286, 33473, 33660, 33847, 34034, 34221, 34408, 34595, 34782, 34969, 35156, 35343, 35530, 35717, 35904, 36091, 36278, 36465, 36652, 36839, 37026, 37213, 37400, 37587, 37774, 37961, 38148, 38335, 38522, 38709, 38896, 39083, 39270, 39457, 39644, 39831, 40018, 40205, 40392, 40579, 40766, 40953, 41140, 41327, 41514, 41701, 41888, 42075, 42262, 42449, 42636, 42823, 43010, 43197, 43384, 43571, 43758, 43945, 44132, 44319, 44506, 44693, 44880, 45067, 45254, 45441, 45628, 45815, 46002, 46189, 46376, 46563, 46750, 46937, 47124, 47311, 47498, 47685, 
0, 188, 376, 564, 752, 940, 1128, 1316, 1504, 1692, 1880, 2068, 2256, 2444, 2632, 2820, 3008, 3196, 3384, 3572, 3760, 3948, 4136, 4324, 4512, 4700, 4888, 5076, 5264, 5452, 5640, 5828, 6016, 6204, 6392, 6580, 6768, 6956, 7144, 7332, 7520, 7708, 7896, 8084, 8272, 8460, 8648, 8836, 9024, 9212, 9400, 9588, 9776, 9964, 10152, 10340, 10528, 10716, 10904, 11092, 11280, 11468, 11656, 11844, 12032, 12220, 12408, 12596, 12784, 12972, 13160, 13348, 13536, 13724, 13912, 14100, 14288, 14476, 14664, 14852, 15040, 15228, 15416, 15604, 15792, 15980, 16168, 16356, 16544, 16732, 16920, 17108, 17296, 17484, 17672, 17860, 18048, 18236, 18424, 18612, 18800, 18988, 19176, 19364, 19552, 19740, 19928, 20116, 20304, 20492, 20680, 20868, 21056, 21244, 21432, 21620, 21808, 21996, 22184, 22372, 22560, 22748, 22936, 23124, 23312, 23500, 23688, 23876, 24064, 24252, 24440, 24628, 24816, 25004, 25192, 25380, 25568, 25756, 25944, 26132, 26320, 26508, 26696, 26884, 27072, 27260, 27448, 27636, 27824, 28012, 28200, 28388, 28576, 28764, 28952, 29140, 29328, 29516, 29704, 29892, 30080, 30268, 30456, 30644, 30832, 31020, 31208, 31396, 31584, 31772, 31960, 32148, 32336, 32524, 32712, 32900, 33088, 33276, 33464, 33652, 33840, 34028, 34216, 34404, 34592, 34780, 34968, 35156, 35344, 35532, 35720, 35908, 36096, 36284, 36472, 36660, 36848, 37036, 37224, 37412, 37600, 37788, 37976, 38164, 38352, 38540, 38728, 38916, 39104, 39292, 39480, 39668, 39856, 40044, 40232, 40420, 40608, 40796, 40984, 41172, 41360, 41548, 41736, 41924, 42112, 42300, 42488, 42676, 42864, 43052, 43240, 43428, 43616, 43804, 43992, 44180, 44368, 44556, 44744, 44932, 45120, 45308, 45496, 45684, 45872, 46060, 46248, 46436, 46624, 46812, 47000, 47188, 47376, 47564, 47752, 47940, 
0, 189, 378, 567, 756, 945, 1134, 1323, 1512, 1701, 1890, 2079, 2268, 2457, 2646, 2835, 3024, 3213, 3402, 3591, 3780, 3969, 4158, 4347, 4536, 4725, 4914, 5103, 5292, 5481, 5670, 5859, 6048, 6237, 6426, 6615, 6804, 6993, 7182, 7371, 7560, 7749, 7938, 8127, 8316, 8505, 8694, 8883, 9072, 9261, 9450, 9639, 9828, 10017, 10206, 10395, 10584, 10773, 10962, 11151, 11340, 11529, 11718, 11907, 12096, 12285, 12474, 12663, 12852, 13041, 13230, 13419, 13608, 13797, 13986, 14175, 14364, 14553, 14742, 14931, 15120, 15309, 15498, 15687, 15876, 16065, 16254, 16443, 16632, 16821, 17010, 17199, 17388, 17577, 17766, 17955, 18144, 18333, 18522, 18711, 18900, 19089, 19278, 19467, 19656, 19845, 20034, 20223, 20412, 20601, 20790, 20979, 21168, 21357, 21546, 21735, 21924, 22113, 22302, 22491, 22680, 22869, 23058, 23247, 23436, 23625, 23814, 24003, 24192, 24381, 24570, 24759, 24948, 25137, 25326, 25515, 25704, 25893, 26082, 26271, 26460, 26649, 26838, 27027, 27216, 27405, 27594, 27783, 27972, 28161, 28350, 28539, 28728, 28917, 29106, 29295, 29484, 29673, 29862, 30051, 30240, 30429, 30618, 30807, 30996, 31185, 31374, 31563, 31752, 31941, 32130, 32319, 32508, 32697, 32886, 33075, 33264, 33453, 33642, 33831, 34020, 34209, 34398, 34587, 34776, 34965, 35154, 35343, 35532, 35721, 35910, 36099, 36288, 36477, 36666, 36855, 37044, 37233, 37422, 37611, 37800, 37989, 38178, 38367, 38556, 38745, 38934, 39123, 39312, 39501, 39690, 39879, 40068, 40257, 40446, 40635, 40824, 41013, 41202, 41391, 41580, 41769, 41958, 42147, 42336, 42525, 42714, 42903, 43092, 43281, 43470, 43659, 43848, 44037, 44226, 44415, 44604, 44793, 44982, 45171, 45360, 45549, 45738, 45927, 46116, 46305, 46494, 46683, 46872, 47061, 47250, 47439, 47628, 47817, 48006, 48195, 
0, 190, 380, 570, 760, 950, 1140, 1330, 1520, 1710, 1900, 2090, 2280, 2470, 2660, 2850, 3040, 3230, 3420, 3610, 3800, 3990, 4180, 4370, 4560, 4750, 4940, 5130, 5320, 5510, 5700, 5890, 6080, 6270, 6460, 6650, 6840, 7030, 7220, 7410, 7600, 7790, 7980, 8170, 8360, 8550, 8740, 8930, 9120, 9310, 9500, 9690, 9880, 10070, 10260, 10450, 10640, 10830, 11020, 11210, 11400, 11590, 11780, 11970, 12160, 12350, 12540, 12730, 12920, 13110, 13300, 13490, 13680, 13870, 14060, 14250, 14440, 14630, 14820, 15010, 15200, 15390, 15580, 15770, 15960, 16150, 16340, 16530, 16720, 16910, 17100, 17290, 17480, 17670, 17860, 18050, 18240, 18430, 18620, 18810, 19000, 19190, 19380, 19570, 19760, 19950, 20140, 20330, 20520, 20710, 20900, 21090, 21280, 21470, 21660, 21850, 22040, 22230, 22420, 22610, 22800, 22990, 23180, 23370, 23560, 23750, 23940, 24130, 24320, 24510, 24700, 24890, 25080, 25270, 25460, 25650, 25840, 26030, 26220, 26410, 26600, 26790, 26980, 27170, 27360, 27550, 27740, 27930, 28120, 28310, 28500, 28690, 28880, 29070, 29260, 29450, 29640, 29830, 30020, 30210, 30400, 30590, 30780, 30970, 31160, 31350, 31540, 31730, 31920, 32110, 32300, 32490, 32680, 32870, 33060, 33250, 33440, 33630, 33820, 34010, 34200, 34390, 34580, 34770, 34960, 35150, 35340, 35530, 35720, 35910, 36100, 36290, 36480, 36670, 36860, 37050, 37240, 37430, 37620, 37810, 38000, 38190, 38380, 38570, 38760, 38950, 39140, 39330, 39520, 39710, 39900, 40090, 40280, 40470, 40660, 40850, 41040, 41230, 41420, 41610, 41800, 41990, 42180, 42370, 42560, 42750, 42940, 43130, 43320, 43510, 43700, 43890, 44080, 44270, 44460, 44650, 44840, 45030, 45220, 45410, 45600, 45790, 45980, 46170, 46360, 46550, 46740, 46930, 47120, 47310, 47500, 47690, 47880, 48070, 48260, 48450, 
0, 191, 382, 573, 764, 955, 1146, 1337, 1528, 1719, 1910, 2101, 2292, 2483, 2674, 2865, 3056, 3247, 3438, 3629, 3820, 4011, 4202, 4393, 4584, 4775, 4966, 5157, 5348, 5539, 5730, 5921, 6112, 6303, 6494, 6685, 6876, 7067, 7258, 7449, 7640, 7831, 8022, 8213, 8404, 8595, 8786, 8977, 9168, 9359, 9550, 9741, 9932, 10123, 10314, 10505, 10696, 10887, 11078, 11269, 11460, 11651, 11842, 12033, 12224, 12415, 12606, 12797, 12988, 13179, 13370, 13561, 13752, 13943, 14134, 14325, 14516, 14707, 14898, 15089, 15280, 15471, 15662, 15853, 16044, 16235, 16426, 16617, 16808, 16999, 17190, 17381, 17572, 17763, 17954, 18145, 18336, 18527, 18718, 18909, 19100, 19291, 19482, 19673, 19864, 20055, 20246, 20437, 20628, 20819, 21010, 21201, 21392, 21583, 21774, 21965, 22156, 22347, 22538, 22729, 22920, 23111, 23302, 23493, 23684, 23875, 24066, 24257, 24448, 24639, 24830, 25021, 25212, 25403, 25594, 25785, 25976, 26167, 26358, 26549, 26740, 26931, 27122, 27313, 27504, 27695, 27886, 28077, 28268, 28459, 28650, 28841, 29032, 29223, 29414, 29605, 29796, 29987, 30178, 30369, 30560, 30751, 30942, 31133, 31324, 31515, 31706, 31897, 32088, 32279, 32470, 32661, 32852, 33043, 33234, 33425, 33616, 33807, 33998, 34189, 34380, 34571, 34762, 34953, 35144, 35335, 35526, 35717, 35908, 36099, 36290, 36481, 36672, 36863, 37054, 37245, 37436, 37627, 37818, 38009, 38200, 38391, 38582, 38773, 38964, 39155, 39346, 39537, 39728, 39919, 40110, 40301, 40492, 40683, 40874, 41065, 41256, 41447, 41638, 41829, 42020, 42211, 42402, 42593, 42784, 42975, 43166, 43357, 43548, 43739, 43930, 44121, 44312, 44503, 44694, 44885, 45076, 45267, 45458, 45649, 45840, 46031, 46222, 46413, 46604, 46795, 46986, 47177, 47368, 47559, 47750, 47941, 48132, 48323, 48514, 48705, 
0, 192, 384, 576, 768, 960, 1152, 1344, 1536, 1728, 1920, 2112, 2304, 2496, 2688, 2880, 3072, 3264, 3456, 3648, 3840, 4032, 4224, 4416, 4608, 4800, 4992, 5184, 5376, 5568, 5760, 5952, 6144, 6336, 6528, 6720, 6912, 7104, 7296, 7488, 7680, 7872, 8064, 8256, 8448, 8640, 8832, 9024, 9216, 9408, 9600, 9792, 9984, 10176, 10368, 10560, 10752, 10944, 11136, 11328, 11520, 11712, 11904, 12096, 12288, 12480, 12672, 12864, 13056, 13248, 13440, 13632, 13824, 14016, 14208, 14400, 14592, 14784, 14976, 15168, 15360, 15552, 15744, 15936, 16128, 16320, 16512, 16704, 16896, 17088, 17280, 17472, 17664, 17856, 18048, 18240, 18432, 18624, 18816, 19008, 19200, 19392, 19584, 19776, 19968, 20160, 20352, 20544, 20736, 20928, 21120, 21312, 21504, 21696, 21888, 22080, 22272, 22464, 22656, 22848, 23040, 23232, 23424, 23616, 23808, 24000, 24192, 24384, 24576, 24768, 24960, 25152, 25344, 25536, 25728, 25920, 26112, 26304, 26496, 26688, 26880, 27072, 27264, 27456, 27648, 27840, 28032, 28224, 28416, 28608, 28800, 28992, 29184, 29376, 29568, 29760, 29952, 30144, 30336, 30528, 30720, 30912, 31104, 31296, 31488, 31680, 31872, 32064, 32256, 32448, 32640, 32832, 33024, 33216, 33408, 33600, 33792, 33984, 34176, 34368, 34560, 34752, 34944, 35136, 35328, 35520, 35712, 35904, 36096, 36288, 36480, 36672, 36864, 37056, 37248, 37440, 37632, 37824, 38016, 38208, 38400, 38592, 38784, 38976, 39168, 39360, 39552, 39744, 39936, 40128, 40320, 40512, 40704, 40896, 41088, 41280, 41472, 41664, 41856, 42048, 42240, 42432, 42624, 42816, 43008, 43200, 43392, 43584, 43776, 43968, 44160, 44352, 44544, 44736, 44928, 45120, 45312, 45504, 45696, 45888, 46080, 46272, 46464, 46656, 46848, 47040, 47232, 47424, 47616, 47808, 48000, 48192, 48384, 48576, 48768, 48960, 
0, 193, 386, 579, 772, 965, 1158, 1351, 1544, 1737, 1930, 2123, 2316, 2509, 2702, 2895, 3088, 3281, 3474, 3667, 3860, 4053, 4246, 4439, 4632, 4825, 5018, 5211, 5404, 5597, 5790, 5983, 6176, 6369, 6562, 6755, 6948, 7141, 7334, 7527, 7720, 7913, 8106, 8299, 8492, 8685, 8878, 9071, 9264, 9457, 9650, 9843, 10036, 10229, 10422, 10615, 10808, 11001, 11194, 11387, 11580, 11773, 11966, 12159, 12352, 12545, 12738, 12931, 13124, 13317, 13510, 13703, 13896, 14089, 14282, 14475, 14668, 14861, 15054, 15247, 15440, 15633, 15826, 16019, 16212, 16405, 16598, 16791, 16984, 17177, 17370, 17563, 17756, 17949, 18142, 18335, 18528, 18721, 18914, 19107, 19300, 19493, 19686, 19879, 20072, 20265, 20458, 20651, 20844, 21037, 21230, 21423, 21616, 21809, 22002, 22195, 22388, 22581, 22774, 22967, 23160, 23353, 23546, 23739, 23932, 24125, 24318, 24511, 24704, 24897, 25090, 25283, 25476, 25669, 25862, 26055, 26248, 26441, 26634, 26827, 27020, 27213, 27406, 27599, 27792, 27985, 28178, 28371, 28564, 28757, 28950, 29143, 29336, 29529, 29722, 29915, 30108, 30301, 30494, 30687, 30880, 31073, 31266, 31459, 31652, 31845, 32038, 32231, 32424, 32617, 32810, 33003, 33196, 33389, 33582, 33775, 33968, 34161, 34354, 34547, 34740, 34933, 35126, 35319, 35512, 35705, 35898, 36091, 36284, 36477, 36670, 36863, 37056, 37249, 37442, 37635, 37828, 38021, 38214, 38407, 38600, 38793, 38986, 39179, 39372, 39565, 39758, 39951, 40144, 40337, 40530, 40723, 40916, 41109, 41302, 41495, 41688, 41881, 42074, 42267, 42460, 42653, 42846, 43039, 43232, 43425, 43618, 43811, 44004, 44197, 44390, 44583, 44776, 44969, 45162, 45355, 45548, 45741, 45934, 46127, 46320, 46513, 46706, 46899, 47092, 47285, 47478, 47671, 47864, 48057, 48250, 48443, 48636, 48829, 49022, 49215, 
0, 194, 388, 582, 776, 970, 1164, 1358, 1552, 1746, 1940, 2134, 2328, 2522, 2716, 2910, 3104, 3298, 3492, 3686, 3880, 4074, 4268, 4462, 4656, 4850, 5044, 5238, 5432, 5626, 5820, 6014, 6208, 6402, 6596, 6790, 6984, 7178, 7372, 7566, 7760, 7954, 8148, 8342, 8536, 8730, 8924, 9118, 9312, 9506, 9700, 9894, 10088, 10282, 10476, 10670, 10864, 11058, 11252, 11446, 11640, 11834, 12028, 12222, 12416, 12610, 12804, 12998, 13192, 13386, 13580, 13774, 13968, 14162, 14356, 14550, 14744, 14938, 15132, 15326, 15520, 15714, 15908, 16102, 16296, 16490, 16684, 16878, 17072, 17266, 17460, 17654, 17848, 18042, 18236, 18430, 18624, 18818, 19012, 19206, 19400, 19594, 19788, 19982, 20176, 20370, 20564, 20758, 20952, 21146, 21340, 21534, 21728, 21922, 22116, 22310, 22504, 22698, 22892, 23086, 23280, 23474, 23668, 23862, 24056, 24250, 24444, 24638, 24832, 25026, 25220, 25414, 25608, 25802, 25996, 26190, 26384, 26578, 26772, 26966, 27160, 27354, 27548, 27742, 27936, 28130, 28324, 28518, 28712, 28906, 29100, 29294, 29488, 29682, 29876, 30070, 30264, 30458, 30652, 30846, 31040, 31234, 31428, 31622, 31816, 32010, 32204, 32398, 32592, 32786, 32980, 33174, 33368, 33562, 33756, 33950, 34144, 34338, 34532, 34726, 34920, 35114, 35308, 35502, 35696, 35890, 36084, 36278, 36472, 36666, 36860, 37054, 37248, 37442, 37636, 37830, 38024, 38218, 38412, 38606, 38800, 38994, 39188, 39382, 39576, 39770, 39964, 40158, 40352, 40546, 40740, 40934, 41128, 41322, 41516, 41710, 41904, 42098, 42292, 42486, 42680, 42874, 43068, 43262, 43456, 43650, 43844, 44038, 44232, 44426, 44620, 44814, 45008, 45202, 45396, 45590, 45784, 45978, 46172, 46366, 46560, 46754, 46948, 47142, 47336, 47530, 47724, 47918, 48112, 48306, 48500, 48694, 48888, 49082, 49276, 49470, 
0, 195, 390, 585, 780, 975, 1170, 1365, 1560, 1755, 1950, 2145, 2340, 2535, 2730, 2925, 3120, 3315, 3510, 3705, 3900, 4095, 4290, 4485, 4680, 4875, 5070, 5265, 5460, 5655, 5850, 6045, 6240, 6435, 6630, 6825, 7020, 7215, 7410, 7605, 7800, 7995, 8190, 8385, 8580, 8775, 8970, 9165, 9360, 9555, 9750, 9945, 10140, 10335, 10530, 10725, 10920, 11115, 11310, 11505, 11700, 11895, 12090, 12285, 12480, 12675, 12870, 13065, 13260, 13455, 13650, 13845, 14040, 14235, 14430, 14625, 14820, 15015, 15210, 15405, 15600, 15795, 15990, 16185, 16380, 16575, 16770, 16965, 17160, 17355, 17550, 17745, 17940, 18135, 18330, 18525, 18720, 18915, 19110, 19305, 19500, 19695, 19890, 20085, 20280, 20475, 20670, 20865, 21060, 21255, 21450, 21645, 21840, 22035, 22230, 22425, 22620, 22815, 23010, 23205, 23400, 23595, 23790, 23985, 24180, 24375, 24570, 24765, 24960, 25155, 25350, 25545, 25740, 25935, 26130, 26325, 26520, 26715, 26910, 27105, 27300, 27495, 27690, 27885, 28080, 28275, 28470, 28665, 28860, 29055, 29250, 29445, 29640, 29835, 30030, 30225, 30420, 30615, 30810, 31005, 31200, 31395, 31590, 31785, 31980, 32175, 32370, 32565, 32760, 32955, 33150, 33345, 33540, 33735, 33930, 34125, 34320, 34515, 34710, 34905, 35100, 35295, 35490, 35685, 35880, 36075, 36270, 36465, 36660, 36855, 37050, 37245, 37440, 37635, 37830, 38025, 38220, 38415, 38610, 38805, 39000, 39195, 39390, 39585, 39780, 39975, 40170, 40365, 40560, 40755, 40950, 41145, 41340, 41535, 41730, 41925, 42120, 42315, 42510, 42705, 42900, 43095, 43290, 43485, 43680, 43875, 44070, 44265, 44460, 44655, 44850, 45045, 45240, 45435, 45630, 45825, 46020, 46215, 46410, 46605, 46800, 46995, 47190, 47385, 47580, 47775, 47970, 48165, 48360, 48555, 48750, 48945, 49140, 49335, 49530, 49725, 
0, 196, 392, 588, 784, 980, 1176, 1372, 1568, 1764, 1960, 2156, 2352, 2548, 2744, 2940, 3136, 3332, 3528, 3724, 3920, 4116, 4312, 4508, 4704, 4900, 5096, 5292, 5488, 5684, 5880, 6076, 6272, 6468, 6664, 6860, 7056, 7252, 7448, 7644, 7840, 8036, 8232, 8428, 8624, 8820, 9016, 9212, 9408, 9604, 9800, 9996, 10192, 10388, 10584, 10780, 10976, 11172, 11368, 11564, 11760, 11956, 12152, 12348, 12544, 12740, 12936, 13132, 13328, 13524, 13720, 13916, 14112, 14308, 14504, 14700, 14896, 15092, 15288, 15484, 15680, 15876, 16072, 16268, 16464, 16660, 16856, 17052, 17248, 17444, 17640, 17836, 18032, 18228, 18424, 18620, 18816, 19012, 19208, 19404, 19600, 19796, 19992, 20188, 20384, 20580, 20776, 20972, 21168, 21364, 21560, 21756, 21952, 22148, 22344, 22540, 22736, 22932, 23128, 23324, 23520, 23716, 23912, 24108, 24304, 24500, 24696, 24892, 25088, 25284, 25480, 25676, 25872, 26068, 26264, 26460, 26656, 26852, 27048, 27244, 27440, 27636, 27832, 28028, 28224, 28420, 28616, 28812, 29008, 29204, 29400, 29596, 29792, 29988, 30184, 30380, 30576, 30772, 30968, 31164, 31360, 31556, 31752, 31948, 32144, 32340, 32536, 32732, 32928, 33124, 33320, 33516, 33712, 33908, 34104, 34300, 34496, 34692, 34888, 35084, 35280, 35476, 35672, 35868, 36064, 36260, 36456, 36652, 36848, 37044, 37240, 37436, 37632, 37828, 38024, 38220, 38416, 38612, 38808, 39004, 39200, 39396, 39592, 39788, 39984, 40180, 40376, 40572, 40768, 40964, 41160, 41356, 41552, 41748, 41944, 42140, 42336, 42532, 42728, 42924, 43120, 43316, 43512, 43708, 43904, 44100, 44296, 44492, 44688, 44884, 45080, 45276, 45472, 45668, 45864, 46060, 46256, 46452, 46648, 46844, 47040, 47236, 47432, 47628, 47824, 48020, 48216, 48412, 48608, 48804, 49000, 49196, 49392, 49588, 49784, 49980, 
0, 197, 394, 591, 788, 985, 1182, 1379, 1576, 1773, 1970, 2167, 2364, 2561, 2758, 2955, 3152, 3349, 3546, 3743, 3940, 4137, 4334, 4531, 4728, 4925, 5122, 5319, 5516, 5713, 5910, 6107, 6304, 6501, 6698, 6895, 7092, 7289, 7486, 7683, 7880, 8077, 8274, 8471, 8668, 8865, 9062, 9259, 9456, 9653, 9850, 10047, 10244, 10441, 10638, 10835, 11032, 11229, 11426, 11623, 11820, 12017, 12214, 12411, 12608, 12805, 13002, 13199, 13396, 13593, 13790, 13987, 14184, 14381, 14578, 14775, 14972, 15169, 15366, 15563, 15760, 15957, 16154, 16351, 16548, 16745, 16942, 17139, 17336, 17533, 17730, 17927, 18124, 18321, 18518, 18715, 18912, 19109, 19306, 19503, 19700, 19897, 20094, 20291, 20488, 20685, 20882, 21079, 21276, 21473, 21670, 21867, 22064, 22261, 22458, 22655, 22852, 23049, 23246, 23443, 23640, 23837, 24034, 24231, 24428, 24625, 24822, 25019, 25216, 25413, 25610, 25807, 26004, 26201, 26398, 26595, 26792, 26989, 27186, 27383, 27580, 27777, 27974, 28171, 28368, 28565, 28762, 28959, 29156, 29353, 29550, 29747, 29944, 30141, 30338, 30535, 30732, 30929, 31126, 31323, 31520, 31717, 31914, 32111, 32308, 32505, 32702, 32899, 33096, 33293, 33490, 33687, 33884, 34081, 34278, 34475, 34672, 34869, 35066, 35263, 35460, 35657, 35854, 36051, 36248, 36445, 36642, 36839, 37036, 37233, 37430, 37627, 37824, 38021, 38218, 38415, 38612, 38809, 39006, 39203, 39400, 39597, 39794, 39991, 40188, 40385, 40582, 40779, 40976, 41173, 41370, 41567, 41764, 41961, 42158, 42355, 42552, 42749, 42946, 43143, 43340, 43537, 43734, 43931, 44128, 44325, 44522, 44719, 44916, 45113, 45310, 45507, 45704, 45901, 46098, 46295, 46492, 46689, 46886, 47083, 47280, 47477, 47674, 47871, 48068, 48265, 48462, 48659, 48856, 49053, 49250, 49447, 49644, 49841, 50038, 50235, 
0, 198, 396, 594, 792, 990, 1188, 1386, 1584, 1782, 1980, 2178, 2376, 2574, 2772, 2970, 3168, 3366, 3564, 3762, 3960, 4158, 4356, 4554, 4752, 4950, 5148, 5346, 5544, 5742, 5940, 6138, 6336, 6534, 6732, 6930, 7128, 7326, 7524, 7722, 7920, 8118, 8316, 8514, 8712, 8910, 9108, 9306, 9504, 9702, 9900, 10098, 10296, 10494, 10692, 10890, 11088, 11286, 11484, 11682, 11880, 12078, 12276, 12474, 12672, 12870, 13068, 13266, 13464, 13662, 13860, 14058, 14256, 14454, 14652, 14850, 15048, 15246, 15444, 15642, 15840, 16038, 16236, 16434, 16632, 16830, 17028, 17226, 17424, 17622, 17820, 18018, 18216, 18414, 18612, 18810, 19008, 19206, 19404, 19602, 19800, 19998, 20196, 20394, 20592, 20790, 20988, 21186, 21384, 21582, 21780, 21978, 22176, 22374, 22572, 22770, 22968, 23166, 23364, 23562, 23760, 23958, 24156, 24354, 24552, 24750, 24948, 25146, 25344, 25542, 25740, 25938, 26136, 26334, 26532, 26730, 26928, 27126, 27324, 27522, 27720, 27918, 28116, 28314, 28512, 28710, 28908, 29106, 29304, 29502, 29700, 29898, 30096, 30294, 30492, 30690, 30888, 31086, 31284, 31482, 31680, 31878, 32076, 32274, 32472, 32670, 32868, 33066, 33264, 33462, 33660, 33858, 34056, 34254, 34452, 34650, 34848, 35046, 35244, 35442, 35640, 35838, 36036, 36234, 36432, 36630, 36828, 37026, 37224, 37422, 37620, 37818, 38016, 38214, 38412, 38610, 38808, 39006, 39204, 39402, 39600, 39798, 39996, 40194, 40392, 40590, 40788, 40986, 41184, 41382, 41580, 41778, 41976, 42174, 42372, 42570, 42768, 42966, 43164, 43362, 43560, 43758, 43956, 44154, 44352, 44550, 44748, 44946, 45144, 45342, 45540, 45738, 45936, 46134, 46332, 46530, 46728, 46926, 47124, 47322, 47520, 47718, 47916, 48114, 48312, 48510, 48708, 48906, 49104, 49302, 49500, 49698, 49896, 50094, 50292, 50490, 
0, 199, 398, 597, 796, 995, 1194, 1393, 1592, 1791, 1990, 2189, 2388, 2587, 2786, 2985, 3184, 3383, 3582, 3781, 3980, 4179, 4378, 4577, 4776, 4975, 5174, 5373, 5572, 5771, 5970, 6169, 6368, 6567, 6766, 6965, 7164, 7363, 7562, 7761, 7960, 8159, 8358, 8557, 8756, 8955, 9154, 9353, 9552, 9751, 9950, 10149, 10348, 10547, 10746, 10945, 11144, 11343, 11542, 11741, 11940, 12139, 12338, 12537, 12736, 12935, 13134, 13333, 13532, 13731, 13930, 14129, 14328, 14527, 14726, 14925, 15124, 15323, 15522, 15721, 15920, 16119, 16318, 16517, 16716, 16915, 17114, 17313, 17512, 17711, 17910, 18109, 18308, 18507, 18706, 18905, 19104, 19303, 19502, 19701, 19900, 20099, 20298, 20497, 20696, 20895, 21094, 21293, 21492, 21691, 21890, 22089, 22288, 22487, 22686, 22885, 23084, 23283, 23482, 23681, 23880, 24079, 24278, 24477, 24676, 24875, 25074, 25273, 25472, 25671, 25870, 26069, 26268, 26467, 26666, 26865, 27064, 27263, 27462, 27661, 27860, 28059, 28258, 28457, 28656, 28855, 29054, 29253, 29452, 29651, 29850, 30049, 30248, 30447, 30646, 30845, 31044, 31243, 31442, 31641, 31840, 32039, 32238, 32437, 32636, 32835, 33034, 33233, 33432, 33631, 33830, 34029, 34228, 34427, 34626, 34825, 35024, 35223, 35422, 35621, 35820, 36019, 36218, 36417, 36616, 36815, 37014, 37213, 37412, 37611, 37810, 38009, 38208, 38407, 38606, 38805, 39004, 39203, 39402, 39601, 39800, 39999, 40198, 40397, 40596, 40795, 40994, 41193, 41392, 41591, 41790, 41989, 42188, 42387, 42586, 42785, 42984, 43183, 43382, 43581, 43780, 43979, 44178, 44377, 44576, 44775, 44974, 45173, 45372, 45571, 45770, 45969, 46168, 46367, 46566, 46765, 46964, 47163, 47362, 47561, 47760, 47959, 48158, 48357, 48556, 48755, 48954, 49153, 49352, 49551, 49750, 49949, 50148, 50347, 50546, 50745, 
0, 200, 400, 600, 800, 1000, 1200, 1400, 1600, 1800, 2000, 2200, 2400, 2600, 2800, 3000, 3200, 3400, 3600, 3800, 4000, 4200, 4400, 4600, 4800, 5000, 5200, 5400, 5600, 5800, 6000, 6200, 6400, 6600, 6800, 7000, 7200, 7400, 7600, 7800, 8000, 8200, 8400, 8600, 8800, 9000, 9200, 9400, 9600, 9800, 10000, 10200, 10400, 10600, 10800, 11000, 11200, 11400, 11600, 11800, 12000, 12200, 12400, 12600, 12800, 13000, 13200, 13400, 13600, 13800, 14000, 14200, 14400, 14600, 14800, 15000, 15200, 15400, 15600, 15800, 16000, 16200, 16400, 16600, 16800, 17000, 17200, 17400, 17600, 17800, 18000, 18200, 18400, 18600, 18800, 19000, 19200, 19400, 19600, 19800, 20000, 20200, 20400, 20600, 20800, 21000, 21200, 21400, 21600, 21800, 22000, 22200, 22400, 22600, 22800, 23000, 23200, 23400, 23600, 23800, 24000, 24200, 24400, 24600, 24800, 25000, 25200, 25400, 25600, 25800, 26000, 26200, 26400, 26600, 26800, 27000, 27200, 27400, 27600, 27800, 28000, 28200, 28400, 28600, 28800, 29000, 29200, 29400, 29600, 29800, 30000, 30200, 30400, 30600, 30800, 31000, 31200, 31400, 31600, 31800, 32000, 32200, 32400, 32600, 32800, 33000, 33200, 33400, 33600, 33800, 34000, 34200, 34400, 34600, 34800, 35000, 35200, 35400, 35600, 35800, 36000, 36200, 36400, 36600, 36800, 37000, 37200, 37400, 37600, 37800, 38000, 38200, 38400, 38600, 38800, 39000, 39200, 39400, 39600, 39800, 40000, 40200, 40400, 40600, 40800, 41000, 41200, 41400, 41600, 41800, 42000, 42200, 42400, 42600, 42800, 43000, 43200, 43400, 43600, 43800, 44000, 44200, 44400, 44600, 44800, 45000, 45200, 45400, 45600, 45800, 46000, 46200, 46400, 46600, 46800, 47000, 47200, 47400, 47600, 47800, 48000, 48200, 48400, 48600, 48800, 49000, 49200, 49400, 49600, 49800, 50000, 50200, 50400, 50600, 50800, 51000, 
0, 201, 402, 603, 804, 1005, 1206, 1407, 1608, 1809, 2010, 2211, 2412, 2613, 2814, 3015, 3216, 3417, 3618, 3819, 4020, 4221, 4422, 4623, 4824, 5025, 5226, 5427, 5628, 5829, 6030, 6231, 6432, 6633, 6834, 7035, 7236, 7437, 7638, 7839, 8040, 8241, 8442, 8643, 8844, 9045, 9246, 9447, 9648, 9849, 10050, 10251, 10452, 10653, 10854, 11055, 11256, 11457, 11658, 11859, 12060, 12261, 12462, 12663, 12864, 13065, 13266, 13467, 13668, 13869, 14070, 14271, 14472, 14673, 14874, 15075, 15276, 15477, 15678, 15879, 16080, 16281, 16482, 16683, 16884, 17085, 17286, 17487, 17688, 17889, 18090, 18291, 18492, 18693, 18894, 19095, 19296, 19497, 19698, 19899, 20100, 20301, 20502, 20703, 20904, 21105, 21306, 21507, 21708, 21909, 22110, 22311, 22512, 22713, 22914, 23115, 23316, 23517, 23718, 23919, 24120, 24321, 24522, 24723, 24924, 25125, 25326, 25527, 25728, 25929, 26130, 26331, 26532, 26733, 26934, 27135, 27336, 27537, 27738, 27939, 28140, 28341, 28542, 28743, 28944, 29145, 29346, 29547, 29748, 29949, 30150, 30351, 30552, 30753, 30954, 31155, 31356, 31557, 31758, 31959, 32160, 32361, 32562, 32763, 32964, 33165, 33366, 33567, 33768, 33969, 34170, 34371, 34572, 34773, 34974, 35175, 35376, 35577, 35778, 35979, 36180, 36381, 36582, 36783, 36984, 37185, 37386, 37587, 37788, 37989, 38190, 38391, 38592, 38793, 38994, 39195, 39396, 39597, 39798, 39999, 40200, 40401, 40602, 40803, 41004, 41205, 41406, 41607, 41808, 42009, 42210, 42411, 42612, 42813, 43014, 43215, 43416, 43617, 43818, 44019, 44220, 44421, 44622, 44823, 45024, 45225, 45426, 45627, 45828, 46029, 46230, 46431, 46632, 46833, 47034, 47235, 47436, 47637, 47838, 48039, 48240, 48441, 48642, 48843, 49044, 49245, 49446, 49647, 49848, 50049, 50250, 50451, 50652, 50853, 51054, 51255, 
0, 202, 404, 606, 808, 1010, 1212, 1414, 1616, 1818, 2020, 2222, 2424, 2626, 2828, 3030, 3232, 3434, 3636, 3838, 4040, 4242, 4444, 4646, 4848, 5050, 5252, 5454, 5656, 5858, 6060, 6262, 6464, 6666, 6868, 7070, 7272, 7474, 7676, 7878, 8080, 8282, 8484, 8686, 8888, 9090, 9292, 9494, 9696, 9898, 10100, 10302, 10504, 10706, 10908, 11110, 11312, 11514, 11716, 11918, 12120, 12322, 12524, 12726, 12928, 13130, 13332, 13534, 13736, 13938, 14140, 14342, 14544, 14746, 14948, 15150, 15352, 15554, 15756, 15958, 16160, 16362, 16564, 16766, 16968, 17170, 17372, 17574, 17776, 17978, 18180, 18382, 18584, 18786, 18988, 19190, 19392, 19594, 19796, 19998, 20200, 20402, 20604, 20806, 21008, 21210, 21412, 21614, 21816, 22018, 22220, 22422, 22624, 22826, 23028, 23230, 23432, 23634, 23836, 24038, 24240, 24442, 24644, 24846, 25048, 25250, 25452, 25654, 25856, 26058, 26260, 26462, 26664, 26866, 27068, 27270, 27472, 27674, 27876, 28078, 28280, 28482, 28684, 28886, 29088, 29290, 29492, 29694, 29896, 30098, 30300, 30502, 30704, 30906, 31108, 31310, 31512, 31714, 31916, 32118, 32320, 32522, 32724, 32926, 33128, 33330, 33532, 33734, 33936, 34138, 34340, 34542, 34744, 34946, 35148, 35350, 35552, 35754, 35956, 36158, 36360, 36562, 36764, 36966, 37168, 37370, 37572, 37774, 37976, 38178, 38380, 38582, 38784, 38986, 39188, 39390, 39592, 39794, 39996, 40198, 40400, 40602, 40804, 41006, 41208, 41410, 41612, 41814, 42016, 42218, 42420, 42622, 42824, 43026, 43228, 43430, 43632, 43834, 44036, 44238, 44440, 44642, 44844, 45046, 45248, 45450, 45652, 45854, 46056, 46258, 46460, 46662, 46864, 47066, 47268, 47470, 47672, 47874, 48076, 48278, 48480, 48682, 48884, 49086, 49288, 49490, 49692, 49894, 50096, 50298, 50500, 50702, 50904, 51106, 51308, 51510, 
0, 203, 406, 609, 812, 1015, 1218, 1421, 1624, 1827, 2030, 2233, 2436, 2639, 2842, 3045, 3248, 3451, 3654, 3857, 4060, 4263, 4466, 4669, 4872, 5075, 5278, 5481, 5684, 5887, 6090, 6293, 6496, 6699, 6902, 7105, 7308, 7511, 7714, 7917, 8120, 8323, 8526, 8729, 8932, 9135, 9338, 9541, 9744, 9947, 10150, 10353, 10556, 10759, 10962, 11165, 11368, 11571, 11774, 11977, 12180, 12383, 12586, 12789, 12992, 13195, 13398, 13601, 13804, 14007, 14210, 14413, 14616, 14819, 15022, 15225, 15428, 15631, 15834, 16037, 16240, 16443, 16646, 16849, 17052, 17255, 17458, 17661, 17864, 18067, 18270, 18473, 18676, 18879, 19082, 19285, 19488, 19691, 19894, 20097, 20300, 20503, 20706, 20909, 21112, 21315, 21518, 21721, 21924, 22127, 22330, 22533, 22736, 22939, 23142, 23345, 23548, 23751, 23954, 24157, 24360, 24563, 24766, 24969, 25172, 25375, 25578, 25781, 25984, 26187, 26390, 26593, 26796, 26999, 27202, 27405, 27608, 27811, 28014, 28217, 28420, 28623, 28826, 29029, 29232, 29435, 29638, 29841, 30044, 30247, 30450, 30653, 30856, 31059, 31262, 31465, 31668, 31871, 32074, 32277, 32480, 32683, 32886, 33089, 33292, 33495, 33698, 33901, 34104, 34307, 34510, 34713, 34916, 35119, 35322, 35525, 35728, 35931, 36134, 36337, 36540, 36743, 36946, 37149, 37352, 37555, 37758, 37961, 38164, 38367, 38570, 38773, 38976, 39179, 39382, 39585, 39788, 39991, 40194, 40397, 40600, 40803, 41006, 41209, 41412, 41615, 41818, 42021, 42224, 42427, 42630, 42833, 43036, 43239, 43442, 43645, 43848, 44051, 44254, 44457, 44660, 44863, 45066, 45269, 45472, 45675, 45878, 46081, 46284, 46487, 46690, 46893, 47096, 47299, 47502, 47705, 47908, 48111, 48314, 48517, 48720, 48923, 49126, 49329, 49532, 49735, 49938, 50141, 50344, 50547, 50750, 50953, 51156, 51359, 51562, 51765, 
0, 204, 408, 612, 816, 1020, 1224, 1428, 1632, 1836, 2040, 2244, 2448, 2652, 2856, 3060, 3264, 3468, 3672, 3876, 4080, 4284, 4488, 4692, 4896, 5100, 5304, 5508, 5712, 5916, 6120, 6324, 6528, 6732, 6936, 7140, 7344, 7548, 7752, 7956, 8160, 8364, 8568, 8772, 8976, 9180, 9384, 9588, 9792, 9996, 10200, 10404, 10608, 10812, 11016, 11220, 11424, 11628, 11832, 12036, 12240, 12444, 12648, 12852, 13056, 13260, 13464, 13668, 13872, 14076, 14280, 14484, 14688, 14892, 15096, 15300, 15504, 15708, 15912, 16116, 16320, 16524, 16728, 16932, 17136, 17340, 17544, 17748, 17952, 18156, 18360, 18564, 18768, 18972, 19176, 19380, 19584, 19788, 19992, 20196, 20400, 20604, 20808, 21012, 21216, 21420, 21624, 21828, 22032, 22236, 22440, 22644, 22848, 23052, 23256, 23460, 23664, 23868, 24072, 24276, 24480, 24684, 24888, 25092, 25296, 25500, 25704, 25908, 26112, 26316, 26520, 26724, 26928, 27132, 27336, 27540, 27744, 27948, 28152, 28356, 28560, 28764, 28968, 29172, 29376, 29580, 29784, 29988, 30192, 30396, 30600, 30804, 31008, 31212, 31416, 31620, 31824, 32028, 32232, 32436, 32640, 32844, 33048, 33252, 33456, 33660, 33864, 34068, 34272, 34476, 34680, 34884, 35088, 35292, 35496, 35700, 35904, 36108, 36312, 36516, 36720, 36924, 37128, 37332, 37536, 37740, 37944, 38148, 38352, 38556, 38760, 38964, 39168, 39372, 39576, 39780, 39984, 40188, 40392, 40596, 40800, 41004, 41208, 41412, 41616, 41820, 42024, 42228, 42432, 42636, 42840, 43044, 43248, 43452, 43656, 43860, 44064, 44268, 44472, 44676, 44880, 45084, 45288, 45492, 45696, 45900, 46104, 46308, 46512, 46716, 46920, 47124, 47328, 47532, 47736, 47940, 48144, 48348, 48552, 48756, 48960, 49164, 49368, 49572, 49776, 49980, 50184, 50388, 50592, 50796, 51000, 51204, 51408, 51612, 51816, 52020, 
0, 205, 410, 615, 820, 1025, 1230, 1435, 1640, 1845, 2050, 2255, 2460, 2665, 2870, 3075, 3280, 3485, 3690, 3895, 4100, 4305, 4510, 4715, 4920, 5125, 5330, 5535, 5740, 5945, 6150, 6355, 6560, 6765, 6970, 7175, 7380, 7585, 7790, 7995, 8200, 8405, 8610, 8815, 9020, 9225, 9430, 9635, 9840, 10045, 10250, 10455, 10660, 10865, 11070, 11275, 11480, 11685, 11890, 12095, 12300, 12505, 12710, 12915, 13120, 13325, 13530, 13735, 13940, 14145, 14350, 14555, 14760, 14965, 15170, 15375, 15580, 15785, 15990, 16195, 16400, 16605, 16810, 17015, 17220, 17425, 17630, 17835, 18040, 18245, 18450, 18655, 18860, 19065, 19270, 19475, 19680, 19885, 20090, 20295, 20500, 20705, 20910, 21115, 21320, 21525, 21730, 21935, 22140, 22345, 22550, 22755, 22960, 23165, 23370, 23575, 23780, 23985, 24190, 24395, 24600, 24805, 25010, 25215, 25420, 25625, 25830, 26035, 26240, 26445, 26650, 26855, 27060, 27265, 27470, 27675, 27880, 28085, 28290, 28495, 28700, 28905, 29110, 29315, 29520, 29725, 29930, 30135, 30340, 30545, 30750, 30955, 31160, 31365, 31570, 31775, 31980, 32185, 32390, 32595, 32800, 33005, 33210, 33415, 33620, 33825, 34030, 34235, 34440, 34645, 34850, 35055, 35260, 35465, 35670, 35875, 36080, 36285, 36490, 36695, 36900, 37105, 37310, 37515, 37720, 37925, 38130, 38335, 38540, 38745, 38950, 39155, 39360, 39565, 39770, 39975, 40180, 40385, 40590, 40795, 41000, 41205, 41410, 41615, 41820, 42025, 42230, 42435, 42640, 42845, 43050, 43255, 43460, 43665, 43870, 44075, 44280, 44485, 44690, 44895, 45100, 45305, 45510, 45715, 45920, 46125, 46330, 46535, 46740, 46945, 47150, 47355, 47560, 47765, 47970, 48175, 48380, 48585, 48790, 48995, 49200, 49405, 49610, 49815, 50020, 50225, 50430, 50635, 50840, 51045, 51250, 51455, 51660, 51865, 52070, 52275, 
0, 206, 412, 618, 824, 1030, 1236, 1442, 1648, 1854, 2060, 2266, 2472, 2678, 2884, 3090, 3296, 3502, 3708, 3914, 4120, 4326, 4532, 4738, 4944, 5150, 5356, 5562, 5768, 5974, 6180, 6386, 6592, 6798, 7004, 7210, 7416, 7622, 7828, 8034, 8240, 8446, 8652, 8858, 9064, 9270, 9476, 9682, 9888, 10094, 10300, 10506, 10712, 10918, 11124, 11330, 11536, 11742, 11948, 12154, 12360, 12566, 12772, 12978, 13184, 13390, 13596, 13802, 14008, 14214, 14420, 14626, 14832, 15038, 15244, 15450, 15656, 15862, 16068, 16274, 16480, 16686, 16892, 17098, 17304, 17510, 17716, 17922, 18128, 18334, 18540, 18746, 18952, 19158, 19364, 19570, 19776, 19982, 20188, 20394, 20600, 20806, 21012, 21218, 21424, 21630, 21836, 22042, 22248, 22454, 22660, 22866, 23072, 23278, 23484, 23690, 23896, 24102, 24308, 24514, 24720, 24926, 25132, 25338, 25544, 25750, 25956, 26162, 26368, 26574, 26780, 26986, 27192, 27398, 27604, 27810, 28016, 28222, 28428, 28634, 28840, 29046, 29252, 29458, 29664, 29870, 30076, 30282, 30488, 30694, 30900, 31106, 31312, 31518, 31724, 31930, 32136, 32342, 32548, 32754, 32960, 33166, 33372, 33578, 33784, 33990, 34196, 34402, 34608, 34814, 35020, 35226, 35432, 35638, 35844, 36050, 36256, 36462, 36668, 36874, 37080, 37286, 37492, 37698, 37904, 38110, 38316, 38522, 38728, 38934, 39140, 39346, 39552, 39758, 39964, 40170, 40376, 40582, 40788, 40994, 41200, 41406, 41612, 41818, 42024, 42230, 42436, 42642, 42848, 43054, 43260, 43466, 43672, 43878, 44084, 44290, 44496, 44702, 44908, 45114, 45320, 45526, 45732, 45938, 46144, 46350, 46556, 46762, 46968, 47174, 47380, 47586, 47792, 47998, 48204, 48410, 48616, 48822, 49028, 49234, 49440, 49646, 49852, 50058, 50264, 50470, 50676, 50882, 51088, 51294, 51500, 51706, 51912, 52118, 52324, 52530, 
0, 207, 414, 621, 828, 1035, 1242, 1449, 1656, 1863, 2070, 2277, 2484, 2691, 2898, 3105, 3312, 3519, 3726, 3933, 4140, 4347, 4554, 4761, 4968, 5175, 5382, 5589, 5796, 6003, 6210, 6417, 6624, 6831, 7038, 7245, 7452, 7659, 7866, 8073, 8280, 8487, 8694, 8901, 9108, 9315, 9522, 9729, 9936, 10143, 10350, 10557, 10764, 10971, 11178, 11385, 11592, 11799, 12006, 12213, 12420, 12627, 12834, 13041, 13248, 13455, 13662, 13869, 14076, 14283, 14490, 14697, 14904, 15111, 15318, 15525, 15732, 15939, 16146, 16353, 16560, 16767, 16974, 17181, 17388, 17595, 17802, 18009, 18216, 18423, 18630, 18837, 19044, 19251, 19458, 19665, 19872, 20079, 20286, 20493, 20700, 20907, 21114, 21321, 21528, 21735, 21942, 22149, 22356, 22563, 22770, 22977, 23184, 23391, 23598, 23805, 24012, 24219, 24426, 24633, 24840, 25047, 25254, 25461, 25668, 25875, 26082, 26289, 26496, 26703, 26910, 27117, 27324, 27531, 27738, 27945, 28152, 28359, 28566, 28773, 28980, 29187, 29394, 29601, 29808, 30015, 30222, 30429, 30636, 30843, 31050, 31257, 31464, 31671, 31878, 32085, 32292, 32499, 32706, 32913, 33120, 33327, 33534, 33741, 33948, 34155, 34362, 34569, 34776, 34983, 35190, 35397, 35604, 35811, 36018, 36225, 36432, 36639, 36846, 37053, 37260, 37467, 37674, 37881, 38088, 38295, 38502, 38709, 38916, 39123, 39330, 39537, 39744, 39951, 40158, 40365, 40572, 40779, 40986, 41193, 41400, 41607, 41814, 42021, 42228, 42435, 42642, 42849, 43056, 43263, 43470, 43677, 43884, 44091, 44298, 44505, 44712, 44919, 45126, 45333, 45540, 45747, 45954, 46161, 46368, 46575, 46782, 46989, 47196, 47403, 47610, 47817, 48024, 48231, 48438, 48645, 48852, 49059, 49266, 49473, 49680, 49887, 50094, 50301, 50508, 50715, 50922, 51129, 51336, 51543, 51750, 51957, 52164, 52371, 52578, 52785, 
0, 208, 416, 624, 832, 1040, 1248, 1456, 1664, 1872, 2080, 2288, 2496, 2704, 2912, 3120, 3328, 3536, 3744, 3952, 4160, 4368, 4576, 4784, 4992, 5200, 5408, 5616, 5824, 6032, 6240, 6448, 6656, 6864, 7072, 7280, 7488, 7696, 7904, 8112, 8320, 8528, 8736, 8944, 9152, 9360, 9568, 9776, 9984, 10192, 10400, 10608, 10816, 11024, 11232, 11440, 11648, 11856, 12064, 12272, 12480, 12688, 12896, 13104, 13312, 13520, 13728, 13936, 14144, 14352, 14560, 14768, 14976, 15184, 15392, 15600, 15808, 16016, 16224, 16432, 16640, 16848, 17056, 17264, 17472, 17680, 17888, 18096, 18304, 18512, 18720, 18928, 19136, 19344, 19552, 19760, 19968, 20176, 20384, 20592, 20800, 21008, 21216, 21424, 21632, 21840, 22048, 22256, 22464, 22672, 22880, 23088, 23296, 23504, 23712, 23920, 24128, 24336, 24544, 24752, 24960, 25168, 25376, 25584, 25792, 26000, 26208, 26416, 26624, 26832, 27040, 27248, 27456, 27664, 27872, 28080, 28288, 28496, 28704, 28912, 29120, 29328, 29536, 29744, 29952, 30160, 30368, 30576, 30784, 30992, 31200, 31408, 31616, 31824, 32032, 32240, 32448, 32656, 32864, 33072, 33280, 33488, 33696, 33904, 34112, 34320, 34528, 34736, 34944, 35152, 35360, 35568, 35776, 35984, 36192, 36400, 36608, 36816, 37024, 37232, 37440, 37648, 37856, 38064, 38272, 38480, 38688, 38896, 39104, 39312, 39520, 39728, 39936, 40144, 40352, 40560, 40768, 40976, 41184, 41392, 41600, 41808, 42016, 42224, 42432, 42640, 42848, 43056, 43264, 43472, 43680, 43888, 44096, 44304, 44512, 44720, 44928, 45136, 45344, 45552, 45760, 45968, 46176, 46384, 46592, 46800, 47008, 47216, 47424, 47632, 47840, 48048, 48256, 48464, 48672, 48880, 49088, 49296, 49504, 49712, 49920, 50128, 50336, 50544, 50752, 50960, 51168, 51376, 51584, 51792, 52000, 52208, 52416, 52624, 52832, 53040, 
0, 209, 418, 627, 836, 1045, 1254, 1463, 1672, 1881, 2090, 2299, 2508, 2717, 2926, 3135, 3344, 3553, 3762, 3971, 4180, 4389, 4598, 4807, 5016, 5225, 5434, 5643, 5852, 6061, 6270, 6479, 6688, 6897, 7106, 7315, 7524, 7733, 7942, 8151, 8360, 8569, 8778, 8987, 9196, 9405, 9614, 9823, 10032, 10241, 10450, 10659, 10868, 11077, 11286, 11495, 11704, 11913, 12122, 12331, 12540, 12749, 12958, 13167, 13376, 13585, 13794, 14003, 14212, 14421, 14630, 14839, 15048, 15257, 15466, 15675, 15884, 16093, 16302, 16511, 16720, 16929, 17138, 17347, 17556, 17765, 17974, 18183, 18392, 18601, 18810, 19019, 19228, 19437, 19646, 19855, 20064, 20273, 20482, 20691, 20900, 21109, 21318, 21527, 21736, 21945, 22154, 22363, 22572, 22781, 22990, 23199, 23408, 23617, 23826, 24035, 24244, 24453, 24662, 24871, 25080, 25289, 25498, 25707, 25916, 26125, 26334, 26543, 26752, 26961, 27170, 27379, 27588, 27797, 28006, 28215, 28424, 28633, 28842, 29051, 29260, 29469, 29678, 29887, 30096, 30305, 30514, 30723, 30932, 31141, 31350, 31559, 31768, 31977, 32186, 32395, 32604, 32813, 33022, 33231, 33440, 33649, 33858, 34067, 34276, 34485, 34694, 34903, 35112, 35321, 35530, 35739, 35948, 36157, 36366, 36575, 36784, 36993, 37202, 37411, 37620, 37829, 38038, 38247, 38456, 38665, 38874, 39083, 39292, 39501, 39710, 39919, 40128, 40337, 40546, 40755, 40964, 41173, 41382, 41591, 41800, 42009, 42218, 42427, 42636, 42845, 43054, 43263, 43472, 43681, 43890, 44099, 44308, 44517, 44726, 44935, 45144, 45353, 45562, 45771, 45980, 46189, 46398, 46607, 46816, 47025, 47234, 47443, 47652, 47861, 48070, 48279, 48488, 48697, 48906, 49115, 49324, 49533, 49742, 49951, 50160, 50369, 50578, 50787, 50996, 51205, 51414, 51623, 51832, 52041, 52250, 52459, 52668, 52877, 53086, 53295, 
0, 210, 420, 630, 840, 1050, 1260, 1470, 1680, 1890, 2100, 2310, 2520, 2730, 2940, 3150, 3360, 3570, 3780, 3990, 4200, 4410, 4620, 4830, 5040, 5250, 5460, 5670, 5880, 6090, 6300, 6510, 6720, 6930, 7140, 7350, 7560, 7770, 7980, 8190, 8400, 8610, 8820, 9030, 9240, 9450, 9660, 9870, 10080, 10290, 10500, 10710, 10920, 11130, 11340, 11550, 11760, 11970, 12180, 12390, 12600, 12810, 13020, 13230, 13440, 13650, 13860, 14070, 14280, 14490, 14700, 14910, 15120, 15330, 15540, 15750, 15960, 16170, 16380, 16590, 16800, 17010, 17220, 17430, 17640, 17850, 18060, 18270, 18480, 18690, 18900, 19110, 19320, 19530, 19740, 19950, 20160, 20370, 20580, 20790, 21000, 21210, 21420, 21630, 21840, 22050, 22260, 22470, 22680, 22890, 23100, 23310, 23520, 23730, 23940, 24150, 24360, 24570, 24780, 24990, 25200, 25410, 25620, 25830, 26040, 26250, 26460, 26670, 26880, 27090, 27300, 27510, 27720, 27930, 28140, 28350, 28560, 28770, 28980, 29190, 29400, 29610, 29820, 30030, 30240, 30450, 30660, 30870, 31080, 31290, 31500, 31710, 31920, 32130, 32340, 32550, 32760, 32970, 33180, 33390, 33600, 33810, 34020, 34230, 34440, 34650, 34860, 35070, 35280, 35490, 35700, 35910, 36120, 36330, 36540, 36750, 36960, 37170, 37380, 37590, 37800, 38010, 38220, 38430, 38640, 38850, 39060, 39270, 39480, 39690, 39900, 40110, 40320, 40530, 40740, 40950, 41160, 41370, 41580, 41790, 42000, 42210, 42420, 42630, 42840, 43050, 43260, 43470, 43680, 43890, 44100, 44310, 44520, 44730, 44940, 45150, 45360, 45570, 45780, 45990, 46200, 46410, 46620, 46830, 47040, 47250, 47460, 47670, 47880, 48090, 48300, 48510, 48720, 48930, 49140, 49350, 49560, 49770, 49980, 50190, 50400, 50610, 50820, 51030, 51240, 51450, 51660, 51870, 52080, 52290, 52500, 52710, 52920, 53130, 53340, 53550, 
0, 211, 422, 633, 844, 1055, 1266, 1477, 1688, 1899, 2110, 2321, 2532, 2743, 2954, 3165, 3376, 3587, 3798, 4009, 4220, 4431, 4642, 4853, 5064, 5275, 5486, 5697, 5908, 6119, 6330, 6541, 6752, 6963, 7174, 7385, 7596, 7807, 8018, 8229, 8440, 8651, 8862, 9073, 9284, 9495, 9706, 9917, 10128, 10339, 10550, 10761, 10972, 11183, 11394, 11605, 11816, 12027, 12238, 12449, 12660, 12871, 13082, 13293, 13504, 13715, 13926, 14137, 14348, 14559, 14770, 14981, 15192, 15403, 15614, 15825, 16036, 16247, 16458, 16669, 16880, 17091, 17302, 17513, 17724, 17935, 18146, 18357, 18568, 18779, 18990, 19201, 19412, 19623, 19834, 20045, 20256, 20467, 20678, 20889, 21100, 21311, 21522, 21733, 21944, 22155, 22366, 22577, 22788, 22999, 23210, 23421, 23632, 23843, 24054, 24265, 24476, 24687, 24898, 25109, 25320, 25531, 25742, 25953, 26164, 26375, 26586, 26797, 27008, 27219, 27430, 27641, 27852, 28063, 28274, 28485, 28696, 28907, 29118, 29329, 29540, 29751, 29962, 30173, 30384, 30595, 30806, 31017, 31228, 31439, 31650, 31861, 32072, 32283, 32494, 32705, 32916, 33127, 33338, 33549, 33760, 33971, 34182, 34393, 34604, 34815, 35026, 35237, 35448, 35659, 35870, 36081, 36292, 36503, 36714, 36925, 37136, 37347, 37558, 37769, 37980, 38191, 38402, 38613, 38824, 39035, 39246, 39457, 39668, 39879, 40090, 40301, 40512, 40723, 40934, 41145, 41356, 41567, 41778, 41989, 42200, 42411, 42622, 42833, 43044, 43255, 43466, 43677, 43888, 44099, 44310, 44521, 44732, 44943, 45154, 45365, 45576, 45787, 45998, 46209, 46420, 46631, 46842, 47053, 47264, 47475, 47686, 47897, 48108, 48319, 48530, 48741, 48952, 49163, 49374, 49585, 49796, 50007, 50218, 50429, 50640, 50851, 51062, 51273, 51484, 51695, 51906, 52117, 52328, 52539, 52750, 52961, 53172, 53383, 53594, 53805, 
0, 212, 424, 636, 848, 1060, 1272, 1484, 1696, 1908, 2120, 2332, 2544, 2756, 2968, 3180, 3392, 3604, 3816, 4028, 4240, 4452, 4664, 4876, 5088, 5300, 5512, 5724, 5936, 6148, 6360, 6572, 6784, 6996, 7208, 7420, 7632, 7844, 8056, 8268, 8480, 8692, 8904, 9116, 9328, 9540, 9752, 9964, 10176, 10388, 10600, 10812, 11024, 11236, 11448, 11660, 11872, 12084, 12296, 12508, 12720, 12932, 13144, 13356, 13568, 13780, 13992, 14204, 14416, 14628, 14840, 15052, 15264, 15476, 15688, 15900, 16112, 16324, 16536, 16748, 16960, 17172, 17384, 17596, 17808, 18020, 18232, 18444, 18656, 18868, 19080, 19292, 19504, 19716, 19928, 20140, 20352, 20564, 20776, 20988, 21200, 21412, 21624, 21836, 22048, 22260, 22472, 22684, 22896, 23108, 23320, 23532, 23744, 23956, 24168, 24380, 24592, 24804, 25016, 25228, 25440, 25652, 25864, 26076, 26288, 26500, 26712, 26924, 27136, 27348, 27560, 27772, 27984, 28196, 28408, 28620, 28832, 29044, 29256, 29468, 29680, 29892, 30104, 30316, 30528, 30740, 30952, 31164, 31376, 31588, 31800, 32012, 32224, 32436, 32648, 32860, 33072, 33284, 33496, 33708, 33920, 34132, 34344, 34556, 34768, 34980, 35192, 35404, 35616, 35828, 36040, 36252, 36464, 36676, 36888, 37100, 37312, 37524, 37736, 37948, 38160, 38372, 38584, 38796, 39008, 39220, 39432, 39644, 39856, 40068, 40280, 40492, 40704, 40916, 41128, 41340, 41552, 41764, 41976, 42188, 42400, 42612, 42824, 43036, 43248, 43460, 43672, 43884, 44096, 44308, 44520, 44732, 44944, 45156, 45368, 45580, 45792, 46004, 46216, 46428, 46640, 46852, 47064, 47276, 47488, 47700, 47912, 48124, 48336, 48548, 48760, 48972, 49184, 49396, 49608, 49820, 50032, 50244, 50456, 50668, 50880, 51092, 51304, 51516, 51728, 51940, 52152, 52364, 52576, 52788, 53000, 53212, 53424, 53636, 53848, 54060, 
0, 213, 426, 639, 852, 1065, 1278, 1491, 1704, 1917, 2130, 2343, 2556, 2769, 2982, 3195, 3408, 3621, 3834, 4047, 4260, 4473, 4686, 4899, 5112, 5325, 5538, 5751, 5964, 6177, 6390, 6603, 6816, 7029, 7242, 7455, 7668, 7881, 8094, 8307, 8520, 8733, 8946, 9159, 9372, 9585, 9798, 10011, 10224, 10437, 10650, 10863, 11076, 11289, 11502, 11715, 11928, 12141, 12354, 12567, 12780, 12993, 13206, 13419, 13632, 13845, 14058, 14271, 14484, 14697, 14910, 15123, 15336, 15549, 15762, 15975, 16188, 16401, 16614, 16827, 17040, 17253, 17466, 17679, 17892, 18105, 18318, 18531, 18744, 18957, 19170, 19383, 19596, 19809, 20022, 20235, 20448, 20661, 20874, 21087, 21300, 21513, 21726, 21939, 22152, 22365, 22578, 22791, 23004, 23217, 23430, 23643, 23856, 24069, 24282, 24495, 24708, 24921, 25134, 25347, 25560, 25773, 25986, 26199, 26412, 26625, 26838, 27051, 27264, 27477, 27690, 27903, 28116, 28329, 28542, 28755, 28968, 29181, 29394, 29607, 29820, 30033, 30246, 30459, 30672, 30885, 31098, 31311, 31524, 31737, 31950, 32163, 32376, 32589, 32802, 33015, 33228, 33441, 33654, 33867, 34080, 34293, 34506, 34719, 34932, 35145, 35358, 35571, 35784, 35997, 36210, 36423, 36636, 36849, 37062, 37275, 37488, 37701, 37914, 38127, 38340, 38553, 38766, 38979, 39192, 39405, 39618, 39831, 40044, 40257, 40470, 40683, 40896, 41109, 41322, 41535, 41748, 41961, 42174, 42387, 42600, 42813, 43026, 43239, 43452, 43665, 43878, 44091, 44304, 44517, 44730, 44943, 45156, 45369, 45582, 45795, 46008, 46221, 46434, 46647, 46860, 47073, 47286, 47499, 47712, 47925, 48138, 48351, 48564, 48777, 48990, 49203, 49416, 49629, 49842, 50055, 50268, 50481, 50694, 50907, 51120, 51333, 51546, 51759, 51972, 52185, 52398, 52611, 52824, 53037, 53250, 53463, 53676, 53889, 54102, 54315, 
0, 214, 428, 642, 856, 1070, 1284, 1498, 1712, 1926, 2140, 2354, 2568, 2782, 2996, 3210, 3424, 3638, 3852, 4066, 4280, 4494, 4708, 4922, 5136, 5350, 5564, 5778, 5992, 6206, 6420, 6634, 6848, 7062, 7276, 7490, 7704, 7918, 8132, 8346, 8560, 8774, 8988, 9202, 9416, 9630, 9844, 10058, 10272, 10486, 10700, 10914, 11128, 11342, 11556, 11770, 11984, 12198, 12412, 12626, 12840, 13054, 13268, 13482, 13696, 13910, 14124, 14338, 14552, 14766, 14980, 15194, 15408, 15622, 15836, 16050, 16264, 16478, 16692, 16906, 17120, 17334, 17548, 17762, 17976, 18190, 18404, 18618, 18832, 19046, 19260, 19474, 19688, 19902, 20116, 20330, 20544, 20758, 20972, 21186, 21400, 21614, 21828, 22042, 22256, 22470, 22684, 22898, 23112, 23326, 23540, 23754, 23968, 24182, 24396, 24610, 24824, 25038, 25252, 25466, 25680, 25894, 26108, 26322, 26536, 26750, 26964, 27178, 27392, 27606, 27820, 28034, 28248, 28462, 28676, 28890, 29104, 29318, 29532, 29746, 29960, 30174, 30388, 30602, 30816, 31030, 31244, 31458, 31672, 31886, 32100, 32314, 32528, 32742, 32956, 33170, 33384, 33598, 33812, 34026, 34240, 34454, 34668, 34882, 35096, 35310, 35524, 35738, 35952, 36166, 36380, 36594, 36808, 37022, 37236, 37450, 37664, 37878, 38092, 38306, 38520, 38734, 38948, 39162, 39376, 39590, 39804, 40018, 40232, 40446, 40660, 40874, 41088, 41302, 41516, 41730, 41944, 42158, 42372, 42586, 42800, 43014, 43228, 43442, 43656, 43870, 44084, 44298, 44512, 44726, 44940, 45154, 45368, 45582, 45796, 46010, 46224, 46438, 46652, 46866, 47080, 47294, 47508, 47722, 47936, 48150, 48364, 48578, 48792, 49006, 49220, 49434, 49648, 49862, 50076, 50290, 50504, 50718, 50932, 51146, 51360, 51574, 51788, 52002, 52216, 52430, 52644, 52858, 53072, 53286, 53500, 53714, 53928, 54142, 54356, 54570, 
0, 215, 430, 645, 860, 1075, 1290, 1505, 1720, 1935, 2150, 2365, 2580, 2795, 3010, 3225, 3440, 3655, 3870, 4085, 4300, 4515, 4730, 4945, 5160, 5375, 5590, 5805, 6020, 6235, 6450, 6665, 6880, 7095, 7310, 7525, 7740, 7955, 8170, 8385, 8600, 8815, 9030, 9245, 9460, 9675, 9890, 10105, 10320, 10535, 10750, 10965, 11180, 11395, 11610, 11825, 12040, 12255, 12470, 12685, 12900, 13115, 13330, 13545, 13760, 13975, 14190, 14405, 14620, 14835, 15050, 15265, 15480, 15695, 15910, 16125, 16340, 16555, 16770, 16985, 17200, 17415, 17630, 17845, 18060, 18275, 18490, 18705, 18920, 19135, 19350, 19565, 19780, 19995, 20210, 20425, 20640, 20855, 21070, 21285, 21500, 21715, 21930, 22145, 22360, 22575, 22790, 23005, 23220, 23435, 23650, 23865, 24080, 24295, 24510, 24725, 24940, 25155, 25370, 25585, 25800, 26015, 26230, 26445, 26660, 26875, 27090, 27305, 27520, 27735, 27950, 28165, 28380, 28595, 28810, 29025, 29240, 29455, 29670, 29885, 30100, 30315, 30530, 30745, 30960, 31175, 31390, 31605, 31820, 32035, 32250, 32465, 32680, 32895, 33110, 33325, 33540, 33755, 33970, 34185, 34400, 34615, 34830, 35045, 35260, 35475, 35690, 35905, 36120, 36335, 36550, 36765, 36980, 37195, 37410, 37625, 37840, 38055, 38270, 38485, 38700, 38915, 39130, 39345, 39560, 39775, 39990, 40205, 40420, 40635, 40850, 41065, 41280, 41495, 41710, 41925, 42140, 42355, 42570, 42785, 43000, 43215, 43430, 43645, 43860, 44075, 44290, 44505, 44720, 44935, 45150, 45365, 45580, 45795, 46010, 46225, 46440, 46655, 46870, 47085, 47300, 47515, 47730, 47945, 48160, 48375, 48590, 48805, 49020, 49235, 49450, 49665, 49880, 50095, 50310, 50525, 50740, 50955, 51170, 51385, 51600, 51815, 52030, 52245, 52460, 52675, 52890, 53105, 53320, 53535, 53750, 53965, 54180, 54395, 54610, 54825, 
0, 216, 432, 648, 864, 1080, 1296, 1512, 1728, 1944, 2160, 2376, 2592, 2808, 3024, 3240, 3456, 3672, 3888, 4104, 4320, 4536, 4752, 4968, 5184, 5400, 5616, 5832, 6048, 6264, 6480, 6696, 6912, 7128, 7344, 7560, 7776, 7992, 8208, 8424, 8640, 8856, 9072, 9288, 9504, 9720, 9936, 10152, 10368, 10584, 10800, 11016, 11232, 11448, 11664, 11880, 12096, 12312, 12528, 12744, 12960, 13176, 13392, 13608, 13824, 14040, 14256, 14472, 14688, 14904, 15120, 15336, 15552, 15768, 15984, 16200, 16416, 16632, 16848, 17064, 17280, 17496, 17712, 17928, 18144, 18360, 18576, 18792, 19008, 19224, 19440, 19656, 19872, 20088, 20304, 20520, 20736, 20952, 21168, 21384, 21600, 21816, 22032, 22248, 22464, 22680, 22896, 23112, 23328, 23544, 23760, 23976, 24192, 24408, 24624, 24840, 25056, 25272, 25488, 25704, 25920, 26136, 26352, 26568, 26784, 27000, 27216, 27432, 27648, 27864, 28080, 28296, 28512, 28728, 28944, 29160, 29376, 29592, 29808, 30024, 30240, 30456, 30672, 30888, 31104, 31320, 31536, 31752, 31968, 32184, 32400, 32616, 32832, 33048, 33264, 33480, 33696, 33912, 34128, 34344, 34560, 34776, 34992, 35208, 35424, 35640, 35856, 36072, 36288, 36504, 36720, 36936, 37152, 37368, 37584, 37800, 38016, 38232, 38448, 38664, 38880, 39096, 39312, 39528, 39744, 39960, 40176, 40392, 40608, 40824, 41040, 41256, 41472, 41688, 41904, 42120, 42336, 42552, 42768, 42984, 43200, 43416, 43632, 43848, 44064, 44280, 44496, 44712, 44928, 45144, 45360, 45576, 45792, 46008, 46224, 46440, 46656, 46872, 47088, 47304, 47520, 47736, 47952, 48168, 48384, 48600, 48816, 49032, 49248, 49464, 49680, 49896, 50112, 50328, 50544, 50760, 50976, 51192, 51408, 51624, 51840, 52056, 52272, 52488, 52704, 52920, 53136, 53352, 53568, 53784, 54000, 54216, 54432, 54648, 54864, 55080, 
0, 217, 434, 651, 868, 1085, 1302, 1519, 1736, 1953, 2170, 2387, 2604, 2821, 3038, 3255, 3472, 3689, 3906, 4123, 4340, 4557, 4774, 4991, 5208, 5425, 5642, 5859, 6076, 6293, 6510, 6727, 6944, 7161, 7378, 7595, 7812, 8029, 8246, 8463, 8680, 8897, 9114, 9331, 9548, 9765, 9982, 10199, 10416, 10633, 10850, 11067, 11284, 11501, 11718, 11935, 12152, 12369, 12586, 12803, 13020, 13237, 13454, 13671, 13888, 14105, 14322, 14539, 14756, 14973, 15190, 15407, 15624, 15841, 16058, 16275, 16492, 16709, 16926, 17143, 17360, 17577, 17794, 18011, 18228, 18445, 18662, 18879, 19096, 19313, 19530, 19747, 19964, 20181, 20398, 20615, 20832, 21049, 21266, 21483, 21700, 21917, 22134, 22351, 22568, 22785, 23002, 23219, 23436, 23653, 23870, 24087, 24304, 24521, 24738, 24955, 25172, 25389, 25606, 25823, 26040, 26257, 26474, 26691, 26908, 27125, 27342, 27559, 27776, 27993, 28210, 28427, 28644, 28861, 29078, 29295, 29512, 29729, 29946, 30163, 30380, 30597, 30814, 31031, 31248, 31465, 31682, 31899, 32116, 32333, 32550, 32767, 32984, 33201, 33418, 33635, 33852, 34069, 34286, 34503, 34720, 34937, 35154, 35371, 35588, 35805, 36022, 36239, 36456, 36673, 36890, 37107, 37324, 37541, 37758, 37975, 38192, 38409, 38626, 38843, 39060, 39277, 39494, 39711, 39928, 40145, 40362, 40579, 40796, 41013, 41230, 41447, 41664, 41881, 42098, 42315, 42532, 42749, 42966, 43183, 43400, 43617, 43834, 44051, 44268, 44485, 44702, 44919, 45136, 45353, 45570, 45787, 46004, 46221, 46438, 46655, 46872, 47089, 47306, 47523, 47740, 47957, 48174, 48391, 48608, 48825, 49042, 49259, 49476, 49693, 49910, 50127, 50344, 50561, 50778, 50995, 51212, 51429, 51646, 51863, 52080, 52297, 52514, 52731, 52948, 53165, 53382, 53599, 53816, 54033, 54250, 54467, 54684, 54901, 55118, 55335, 
0, 218, 436, 654, 872, 1090, 1308, 1526, 1744, 1962, 2180, 2398, 2616, 2834, 3052, 3270, 3488, 3706, 3924, 4142, 4360, 4578, 4796, 5014, 5232, 5450, 5668, 5886, 6104, 6322, 6540, 6758, 6976, 7194, 7412, 7630, 7848, 8066, 8284, 8502, 8720, 8938, 9156, 9374, 9592, 9810, 10028, 10246, 10464, 10682, 10900, 11118, 11336, 11554, 11772, 11990, 12208, 12426, 12644, 12862, 13080, 13298, 13516, 13734, 13952, 14170, 14388, 14606, 14824, 15042, 15260, 15478, 15696, 15914, 16132, 16350, 16568, 16786, 17004, 17222, 17440, 17658, 17876, 18094, 18312, 18530, 18748, 18966, 19184, 19402, 19620, 19838, 20056, 20274, 20492, 20710, 20928, 21146, 21364, 21582, 21800, 22018, 22236, 22454, 22672, 22890, 23108, 23326, 23544, 23762, 23980, 24198, 24416, 24634, 24852, 25070, 25288, 25506, 25724, 25942, 26160, 26378, 26596, 26814, 27032, 27250, 27468, 27686, 27904, 28122, 28340, 28558, 28776, 28994, 29212, 29430, 29648, 29866, 30084, 30302, 30520, 30738, 30956, 31174, 31392, 31610, 31828, 32046, 32264, 32482, 32700, 32918, 33136, 33354, 33572, 33790, 34008, 34226, 34444, 34662, 34880, 35098, 35316, 35534, 35752, 35970, 36188, 36406, 36624, 36842, 37060, 37278, 37496, 37714, 37932, 38150, 38368, 38586, 38804, 39022, 39240, 39458, 39676, 39894, 40112, 40330, 40548, 40766, 40984, 41202, 41420, 41638, 41856, 42074, 42292, 42510, 42728, 42946, 43164, 43382, 43600, 43818, 44036, 44254, 44472, 44690, 44908, 45126, 45344, 45562, 45780, 45998, 46216, 46434, 46652, 46870, 47088, 47306, 47524, 47742, 47960, 48178, 48396, 48614, 48832, 49050, 49268, 49486, 49704, 49922, 50140, 50358, 50576, 50794, 51012, 51230, 51448, 51666, 51884, 52102, 52320, 52538, 52756, 52974, 53192, 53410, 53628, 53846, 54064, 54282, 54500, 54718, 54936, 55154, 55372, 55590, 
0, 219, 438, 657, 876, 1095, 1314, 1533, 1752, 1971, 2190, 2409, 2628, 2847, 3066, 3285, 3504, 3723, 3942, 4161, 4380, 4599, 4818, 5037, 5256, 5475, 5694, 5913, 6132, 6351, 6570, 6789, 7008, 7227, 7446, 7665, 7884, 8103, 8322, 8541, 8760, 8979, 9198, 9417, 9636, 9855, 10074, 10293, 10512, 10731, 10950, 11169, 11388, 11607, 11826, 12045, 12264, 12483, 12702, 12921, 13140, 13359, 13578, 13797, 14016, 14235, 14454, 14673, 14892, 15111, 15330, 15549, 15768, 15987, 16206, 16425, 16644, 16863, 17082, 17301, 17520, 17739, 17958, 18177, 18396, 18615, 18834, 19053, 19272, 19491, 19710, 19929, 20148, 20367, 20586, 20805, 21024, 21243, 21462, 21681, 21900, 22119, 22338, 22557, 22776, 22995, 23214, 23433, 23652, 23871, 24090, 24309, 24528, 24747, 24966, 25185, 25404, 25623, 25842, 26061, 26280, 26499, 26718, 26937, 27156, 27375, 27594, 27813, 28032, 28251, 28470, 28689, 28908, 29127, 29346, 29565, 29784, 30003, 30222, 30441, 30660, 30879, 31098, 31317, 31536, 31755, 31974, 32193, 32412, 32631, 32850, 33069, 33288, 33507, 33726, 33945, 34164, 34383, 34602, 34821, 35040, 35259, 35478, 35697, 35916, 36135, 36354, 36573, 36792, 37011, 37230, 37449, 37668, 37887, 38106, 38325, 38544, 38763, 38982, 39201, 39420, 39639, 39858, 40077, 40296, 40515, 40734, 40953, 41172, 41391, 41610, 41829, 42048, 42267, 42486, 42705, 42924, 43143, 43362, 43581, 43800, 44019, 44238, 44457, 44676, 44895, 45114, 45333, 45552, 45771, 45990, 46209, 46428, 46647, 46866, 47085, 47304, 47523, 47742, 47961, 48180, 48399, 48618, 48837, 49056, 49275, 49494, 49713, 49932, 50151, 50370, 50589, 50808, 51027, 51246, 51465, 51684, 51903, 52122, 52341, 52560, 52779, 52998, 53217, 53436, 53655, 53874, 54093, 54312, 54531, 54750, 54969, 55188, 55407, 55626, 55845, 
0, 220, 440, 660, 880, 1100, 1320, 1540, 1760, 1980, 2200, 2420, 2640, 2860, 3080, 3300, 3520, 3740, 3960, 4180, 4400, 4620, 4840, 5060, 5280, 5500, 5720, 5940, 6160, 6380, 6600, 6820, 7040, 7260, 7480, 7700, 7920, 8140, 8360, 8580, 8800, 9020, 9240, 9460, 9680, 9900, 10120, 10340, 10560, 10780, 11000, 11220, 11440, 11660, 11880, 12100, 12320, 12540, 12760, 12980, 13200, 13420, 13640, 13860, 14080, 14300, 14520, 14740, 14960, 15180, 15400, 15620, 15840, 16060, 16280, 16500, 16720, 16940, 17160, 17380, 17600, 17820, 18040, 18260, 18480, 18700, 18920, 19140, 19360, 19580, 19800, 20020, 20240, 20460, 20680, 20900, 21120, 21340, 21560, 21780, 22000, 22220, 22440, 22660, 22880, 23100, 23320, 23540, 23760, 23980, 24200, 24420, 24640, 24860, 25080, 25300, 25520, 25740, 25960, 26180, 26400, 26620, 26840, 27060, 27280, 27500, 27720, 27940, 28160, 28380, 28600, 28820, 29040, 29260, 29480, 29700, 29920, 30140, 30360, 30580, 30800, 31020, 31240, 31460, 31680, 31900, 32120, 32340, 32560, 32780, 33000, 33220, 33440, 33660, 33880, 34100, 34320, 34540, 34760, 34980, 35200, 35420, 35640, 35860, 36080, 36300, 36520, 36740, 36960, 37180, 37400, 37620, 37840, 38060, 38280, 38500, 38720, 38940, 39160, 39380, 39600, 39820, 40040, 40260, 40480, 40700, 40920, 41140, 41360, 41580, 41800, 42020, 42240, 42460, 42680, 42900, 43120, 43340, 43560, 43780, 44000, 44220, 44440, 44660, 44880, 45100, 45320, 45540, 45760, 45980, 46200, 46420, 46640, 46860, 47080, 47300, 47520, 47740, 47960, 48180, 48400, 48620, 48840, 49060, 49280, 49500, 49720, 49940, 50160, 50380, 50600, 50820, 51040, 51260, 51480, 51700, 51920, 52140, 52360, 52580, 52800, 53020, 53240, 53460, 53680, 53900, 54120, 54340, 54560, 54780, 55000, 55220, 55440, 55660, 55880, 56100, 
0, 221, 442, 663, 884, 1105, 1326, 1547, 1768, 1989, 2210, 2431, 2652, 2873, 3094, 3315, 3536, 3757, 3978, 4199, 4420, 4641, 4862, 5083, 5304, 5525, 5746, 5967, 6188, 6409, 6630, 6851, 7072, 7293, 7514, 7735, 7956, 8177, 8398, 8619, 8840, 9061, 9282, 9503, 9724, 9945, 10166, 10387, 10608, 10829, 11050, 11271, 11492, 11713, 11934, 12155, 12376, 12597, 12818, 13039, 13260, 13481, 13702, 13923, 14144, 14365, 14586, 14807, 15028, 15249, 15470, 15691, 15912, 16133, 16354, 16575, 16796, 17017, 17238, 17459, 17680, 17901, 18122, 18343, 18564, 18785, 19006, 19227, 19448, 19669, 19890, 20111, 20332, 20553, 20774, 20995, 21216, 21437, 21658, 21879, 22100, 22321, 22542, 22763, 22984, 23205, 23426, 23647, 23868, 24089, 24310, 24531, 24752, 24973, 25194, 25415, 25636, 25857, 26078, 26299, 26520, 26741, 26962, 27183, 27404, 27625, 27846, 28067, 28288, 28509, 28730, 28951, 29172, 29393, 29614, 29835, 30056, 30277, 30498, 30719, 30940, 31161, 31382, 31603, 31824, 32045, 32266, 32487, 32708, 32929, 33150, 33371, 33592, 33813, 34034, 34255, 34476, 34697, 34918, 35139, 35360, 35581, 35802, 36023, 36244, 36465, 36686, 36907, 37128, 37349, 37570, 37791, 38012, 38233, 38454, 38675, 38896, 39117, 39338, 39559, 39780, 40001, 40222, 40443, 40664, 40885, 41106, 41327, 41548, 41769, 41990, 42211, 42432, 42653, 42874, 43095, 43316, 43537, 43758, 43979, 44200, 44421, 44642, 44863, 45084, 45305, 45526, 45747, 45968, 46189, 46410, 46631, 46852, 47073, 47294, 47515, 47736, 47957, 48178, 48399, 48620, 48841, 49062, 49283, 49504, 49725, 49946, 50167, 50388, 50609, 50830, 51051, 51272, 51493, 51714, 51935, 52156, 52377, 52598, 52819, 53040, 53261, 53482, 53703, 53924, 54145, 54366, 54587, 54808, 55029, 55250, 55471, 55692, 55913, 56134, 56355, 
0, 222, 444, 666, 888, 1110, 1332, 1554, 1776, 1998, 2220, 2442, 2664, 2886, 3108, 3330, 3552, 3774, 3996, 4218, 4440, 4662, 4884, 5106, 5328, 5550, 5772, 5994, 6216, 6438, 6660, 6882, 7104, 7326, 7548, 7770, 7992, 8214, 8436, 8658, 8880, 9102, 9324, 9546, 9768, 9990, 10212, 10434, 10656, 10878, 11100, 11322, 11544, 11766, 11988, 12210, 12432, 12654, 12876, 13098, 13320, 13542, 13764, 13986, 14208, 14430, 14652, 14874, 15096, 15318, 15540, 15762, 15984, 16206, 16428, 16650, 16872, 17094, 17316, 17538, 17760, 17982, 18204, 18426, 18648, 18870, 19092, 19314, 19536, 19758, 19980, 20202, 20424, 20646, 20868, 21090, 21312, 21534, 21756, 21978, 22200, 22422, 22644, 22866, 23088, 23310, 23532, 23754, 23976, 24198, 24420, 24642, 24864, 25086, 25308, 25530, 25752, 25974, 26196, 26418, 26640, 26862, 27084, 27306, 27528, 27750, 27972, 28194, 28416, 28638, 28860, 29082, 29304, 29526, 29748, 29970, 30192, 30414, 30636, 30858, 31080, 31302, 31524, 31746, 31968, 32190, 32412, 32634, 32856, 33078, 33300, 33522, 33744, 33966, 34188, 34410, 34632, 34854, 35076, 35298, 35520, 35742, 35964, 36186, 36408, 36630, 36852, 37074, 37296, 37518, 37740, 37962, 38184, 38406, 38628, 38850, 39072, 39294, 39516, 39738, 39960, 40182, 40404, 40626, 40848, 41070, 41292, 41514, 41736, 41958, 42180, 42402, 42624, 42846, 43068, 43290, 43512, 43734, 43956, 44178, 44400, 44622, 44844, 45066, 45288, 45510, 45732, 45954, 46176, 46398, 46620, 46842, 47064, 47286, 47508, 47730, 47952, 48174, 48396, 48618, 48840, 49062, 49284, 49506, 49728, 49950, 50172, 50394, 50616, 50838, 51060, 51282, 51504, 51726, 51948, 52170, 52392, 52614, 52836, 53058, 53280, 53502, 53724, 53946, 54168, 54390, 54612, 54834, 55056, 55278, 55500, 55722, 55944, 56166, 56388, 56610, 
0, 223, 446, 669, 892, 1115, 1338, 1561, 1784, 2007, 2230, 2453, 2676, 2899, 3122, 3345, 3568, 3791, 4014, 4237, 4460, 4683, 4906, 5129, 5352, 5575, 5798, 6021, 6244, 6467, 6690, 6913, 7136, 7359, 7582, 7805, 8028, 8251, 8474, 8697, 8920, 9143, 9366, 9589, 9812, 10035, 10258, 10481, 10704, 10927, 11150, 11373, 11596, 11819, 12042, 12265, 12488, 12711, 12934, 13157, 13380, 13603, 13826, 14049, 14272, 14495, 14718, 14941, 15164, 15387, 15610, 15833, 16056, 16279, 16502, 16725, 16948, 17171, 17394, 17617, 17840, 18063, 18286, 18509, 18732, 18955, 19178, 19401, 19624, 19847, 20070, 20293, 20516, 20739, 20962, 21185, 21408, 21631, 21854, 22077, 22300, 22523, 22746, 22969, 23192, 23415, 23638, 23861, 24084, 24307, 24530, 24753, 24976, 25199, 25422, 25645, 25868, 26091, 26314, 26537, 26760, 26983, 27206, 27429, 27652, 27875, 28098, 28321, 28544, 28767, 28990, 29213, 29436, 29659, 29882, 30105, 30328, 30551, 30774, 30997, 31220, 31443, 31666, 31889, 32112, 32335, 32558, 32781, 33004, 33227, 33450, 33673, 33896, 34119, 34342, 34565, 34788, 35011, 35234, 35457, 35680, 35903, 36126, 36349, 36572, 36795, 37018, 37241, 37464, 37687, 37910, 38133, 38356, 38579, 38802, 39025, 39248, 39471, 39694, 39917, 40140, 40363, 40586, 40809, 41032, 41255, 41478, 41701, 41924, 42147, 42370, 42593, 42816, 43039, 43262, 43485, 43708, 43931, 44154, 44377, 44600, 44823, 45046, 45269, 45492, 45715, 45938, 46161, 46384, 46607, 46830, 47053, 47276, 47499, 47722, 47945, 48168, 48391, 48614, 48837, 49060, 49283, 49506, 49729, 49952, 50175, 50398, 50621, 50844, 51067, 51290, 51513, 51736, 51959, 52182, 52405, 52628, 52851, 53074, 53297, 53520, 53743, 53966, 54189, 54412, 54635, 54858, 55081, 55304, 55527, 55750, 55973, 56196, 56419, 56642, 56865, 
0, 224, 448, 672, 896, 1120, 1344, 1568, 1792, 2016, 2240, 2464, 2688, 2912, 3136, 3360, 3584, 3808, 4032, 4256, 4480, 4704, 4928, 5152, 5376, 5600, 5824, 6048, 6272, 6496, 6720, 6944, 7168, 7392, 7616, 7840, 8064, 8288, 8512, 8736, 8960, 9184, 9408, 9632, 9856, 10080, 10304, 10528, 10752, 10976, 11200, 11424, 11648, 11872, 12096, 12320, 12544, 12768, 12992, 13216, 13440, 13664, 13888, 14112, 14336, 14560, 14784, 15008, 15232, 15456, 15680, 15904, 16128, 16352, 16576, 16800, 17024, 17248, 17472, 17696, 17920, 18144, 18368, 18592, 18816, 19040, 19264, 19488, 19712, 19936, 20160, 20384, 20608, 20832, 21056, 21280, 21504, 21728, 21952, 22176, 22400, 22624, 22848, 23072, 23296, 23520, 23744, 23968, 24192, 24416, 24640, 24864, 25088, 25312, 25536, 25760, 25984, 26208, 26432, 26656, 26880, 27104, 27328, 27552, 27776, 28000, 28224, 28448, 28672, 28896, 29120, 29344, 29568, 29792, 30016, 30240, 30464, 30688, 30912, 31136, 31360, 31584, 31808, 32032, 32256, 32480, 32704, 32928, 33152, 33376, 33600, 33824, 34048, 34272, 34496, 34720, 34944, 35168, 35392, 35616, 35840, 36064, 36288, 36512, 36736, 36960, 37184, 37408, 37632, 37856, 38080, 38304, 38528, 38752, 38976, 39200, 39424, 39648, 39872, 40096, 40320, 40544, 40768, 40992, 41216, 41440, 41664, 41888, 42112, 42336, 42560, 42784, 43008, 43232, 43456, 43680, 43904, 44128, 44352, 44576, 44800, 45024, 45248, 45472, 45696, 45920, 46144, 46368, 46592, 46816, 47040, 47264, 47488, 47712, 47936, 48160, 48384, 48608, 48832, 49056, 49280, 49504, 49728, 49952, 50176, 50400, 50624, 50848, 51072, 51296, 51520, 51744, 51968, 52192, 52416, 52640, 52864, 53088, 53312, 53536, 53760, 53984, 54208, 54432, 54656, 54880, 55104, 55328, 55552, 55776, 56000, 56224, 56448, 56672, 56896, 57120, 
0, 225, 450, 675, 900, 1125, 1350, 1575, 1800, 2025, 2250, 2475, 2700, 2925, 3150, 3375, 3600, 3825, 4050, 4275, 4500, 4725, 4950, 5175, 5400, 5625, 5850, 6075, 6300, 6525, 6750, 6975, 7200, 7425, 7650, 7875, 8100, 8325, 8550, 8775, 9000, 9225, 9450, 9675, 9900, 10125, 10350, 10575, 10800, 11025, 11250, 11475, 11700, 11925, 12150, 12375, 12600, 12825, 13050, 13275, 13500, 13725, 13950, 14175, 14400, 14625, 14850, 15075, 15300, 15525, 15750, 15975, 16200, 16425, 16650, 16875, 17100, 17325, 17550, 17775, 18000, 18225, 18450, 18675, 18900, 19125, 19350, 19575, 19800, 20025, 20250, 20475, 20700, 20925, 21150, 21375, 21600, 21825, 22050, 22275, 22500, 22725, 22950, 23175, 23400, 23625, 23850, 24075, 24300, 24525, 24750, 24975, 25200, 25425, 25650, 25875, 26100, 26325, 26550, 26775, 27000, 27225, 27450, 27675, 27900, 28125, 28350, 28575, 28800, 29025, 29250, 29475, 29700, 29925, 30150, 30375, 30600, 30825, 31050, 31275, 31500, 31725, 31950, 32175, 32400, 32625, 32850, 33075, 33300, 33525, 33750, 33975, 34200, 34425, 34650, 34875, 35100, 35325, 35550, 35775, 36000, 36225, 36450, 36675, 36900, 37125, 37350, 37575, 37800, 38025, 38250, 38475, 38700, 38925, 39150, 39375, 39600, 39825, 40050, 40275, 40500, 40725, 40950, 41175, 41400, 41625, 41850, 42075, 42300, 42525, 42750, 42975, 43200, 43425, 43650, 43875, 44100, 44325, 44550, 44775, 45000, 45225, 45450, 45675, 45900, 46125, 46350, 46575, 46800, 47025, 47250, 47475, 47700, 47925, 48150, 48375, 48600, 48825, 49050, 49275, 49500, 49725, 49950, 50175, 50400, 50625, 50850, 51075, 51300, 51525, 51750, 51975, 52200, 52425, 52650, 52875, 53100, 53325, 53550, 53775, 54000, 54225, 54450, 54675, 54900, 55125, 55350, 55575, 55800, 56025, 56250, 56475, 56700, 56925, 57150, 57375, 
0, 226, 452, 678, 904, 1130, 1356, 1582, 1808, 2034, 2260, 2486, 2712, 2938, 3164, 3390, 3616, 3842, 4068, 4294, 4520, 4746, 4972, 5198, 5424, 5650, 5876, 6102, 6328, 6554, 6780, 7006, 7232, 7458, 7684, 7910, 8136, 8362, 8588, 8814, 9040, 9266, 9492, 9718, 9944, 10170, 10396, 10622, 10848, 11074, 11300, 11526, 11752, 11978, 12204, 12430, 12656, 12882, 13108, 13334, 13560, 13786, 14012, 14238, 14464, 14690, 14916, 15142, 15368, 15594, 15820, 16046, 16272, 16498, 16724, 16950, 17176, 17402, 17628, 17854, 18080, 18306, 18532, 18758, 18984, 19210, 19436, 19662, 19888, 20114, 20340, 20566, 20792, 21018, 21244, 21470, 21696, 21922, 22148, 22374, 22600, 22826, 23052, 23278, 23504, 23730, 23956, 24182, 24408, 24634, 24860, 25086, 25312, 25538, 25764, 25990, 26216, 26442, 26668, 26894, 27120, 27346, 27572, 27798, 28024, 28250, 28476, 28702, 28928, 29154, 29380, 29606, 29832, 30058, 30284, 30510, 30736, 30962, 31188, 31414, 31640, 31866, 32092, 32318, 32544, 32770, 32996, 33222, 33448, 33674, 33900, 34126, 34352, 34578, 34804, 35030, 35256, 35482, 35708, 35934, 36160, 36386, 36612, 36838, 37064, 37290, 37516, 37742, 37968, 38194, 38420, 38646, 38872, 39098, 39324, 39550, 39776, 40002, 40228, 40454, 40680, 40906, 41132, 41358, 41584, 41810, 42036, 42262, 42488, 42714, 42940, 43166, 43392, 43618, 43844, 44070, 44296, 44522, 44748, 44974, 45200, 45426, 45652, 45878, 46104, 46330, 46556, 46782, 47008, 47234, 47460, 47686, 47912, 48138, 48364, 48590, 48816, 49042, 49268, 49494, 49720, 49946, 50172, 50398, 50624, 50850, 51076, 51302, 51528, 51754, 51980, 52206, 52432, 52658, 52884, 53110, 53336, 53562, 53788, 54014, 54240, 54466, 54692, 54918, 55144, 55370, 55596, 55822, 56048, 56274, 56500, 56726, 56952, 57178, 57404, 57630, 
0, 227, 454, 681, 908, 1135, 1362, 1589, 1816, 2043, 2270, 2497, 2724, 2951, 3178, 3405, 3632, 3859, 4086, 4313, 4540, 4767, 4994, 5221, 5448, 5675, 5902, 6129, 6356, 6583, 6810, 7037, 7264, 7491, 7718, 7945, 8172, 8399, 8626, 8853, 9080, 9307, 9534, 9761, 9988, 10215, 10442, 10669, 10896, 11123, 11350, 11577, 11804, 12031, 12258, 12485, 12712, 12939, 13166, 13393, 13620, 13847, 14074, 14301, 14528, 14755, 14982, 15209, 15436, 15663, 15890, 16117, 16344, 16571, 16798, 17025, 17252, 17479, 17706, 17933, 18160, 18387, 18614, 18841, 19068, 19295, 19522, 19749, 19976, 20203, 20430, 20657, 20884, 21111, 21338, 21565, 21792, 22019, 22246, 22473, 22700, 22927, 23154, 23381, 23608, 23835, 24062, 24289, 24516, 24743, 24970, 25197, 25424, 25651, 25878, 26105, 26332, 26559, 26786, 27013, 27240, 27467, 27694, 27921, 28148, 28375, 28602, 28829, 29056, 29283, 29510, 29737, 29964, 30191, 30418, 30645, 30872, 31099, 31326, 31553, 31780, 32007, 32234, 32461, 32688, 32915, 33142, 33369, 33596, 33823, 34050, 34277, 34504, 34731, 34958, 35185, 35412, 35639, 35866, 36093, 36320, 36547, 36774, 37001, 37228, 37455, 37682, 37909, 38136, 38363, 38590, 38817, 39044, 39271, 39498, 39725, 39952, 40179, 40406, 40633, 40860, 41087, 41314, 41541, 41768, 41995, 42222, 42449, 42676, 42903, 43130, 43357, 43584, 43811, 44038, 44265, 44492, 44719, 44946, 45173, 45400, 45627, 45854, 46081, 46308, 46535, 46762, 46989, 47216, 47443, 47670, 47897, 48124, 48351, 48578, 48805, 49032, 49259, 49486, 49713, 49940, 50167, 50394, 50621, 50848, 51075, 51302, 51529, 51756, 51983, 52210, 52437, 52664, 52891, 53118, 53345, 53572, 53799, 54026, 54253, 54480, 54707, 54934, 55161, 55388, 55615, 55842, 56069, 56296, 56523, 56750, 56977, 57204, 57431, 57658, 57885, 
0, 228, 456, 684, 912, 1140, 1368, 1596, 1824, 2052, 2280, 2508, 2736, 2964, 3192, 3420, 3648, 3876, 4104, 4332, 4560, 4788, 5016, 5244, 5472, 5700, 5928, 6156, 6384, 6612, 6840, 7068, 7296, 7524, 7752, 7980, 8208, 8436, 8664, 8892, 9120, 9348, 9576, 9804, 10032, 10260, 10488, 10716, 10944, 11172, 11400, 11628, 11856, 12084, 12312, 12540, 12768, 12996, 13224, 13452, 13680, 13908, 14136, 14364, 14592, 14820, 15048, 15276, 15504, 15732, 15960, 16188, 16416, 16644, 16872, 17100, 17328, 17556, 17784, 18012, 18240, 18468, 18696, 18924, 19152, 19380, 19608, 19836, 20064, 20292, 20520, 20748, 20976, 21204, 21432, 21660, 21888, 22116, 22344, 22572, 22800, 23028, 23256, 23484, 23712, 23940, 24168, 24396, 24624, 24852, 25080, 25308, 25536, 25764, 25992, 26220, 26448, 26676, 26904, 27132, 27360, 27588, 27816, 28044, 28272, 28500, 28728, 28956, 29184, 29412, 29640, 29868, 30096, 30324, 30552, 30780, 31008, 31236, 31464, 31692, 31920, 32148, 32376, 32604, 32832, 33060, 33288, 33516, 33744, 33972, 34200, 34428, 34656, 34884, 35112, 35340, 35568, 35796, 36024, 36252, 36480, 36708, 36936, 37164, 37392, 37620, 37848, 38076, 38304, 38532, 38760, 38988, 39216, 39444, 39672, 39900, 40128, 40356, 40584, 40812, 41040, 41268, 41496, 41724, 41952, 42180, 42408, 42636, 42864, 43092, 43320, 43548, 43776, 44004, 44232, 44460, 44688, 44916, 45144, 45372, 45600, 45828, 46056, 46284, 46512, 46740, 46968, 47196, 47424, 47652, 47880, 48108, 48336, 48564, 48792, 49020, 49248, 49476, 49704, 49932, 50160, 50388, 50616, 50844, 51072, 51300, 51528, 51756, 51984, 52212, 52440, 52668, 52896, 53124, 53352, 53580, 53808, 54036, 54264, 54492, 54720, 54948, 55176, 55404, 55632, 55860, 56088, 56316, 56544, 56772, 57000, 57228, 57456, 57684, 57912, 58140, 
0, 229, 458, 687, 916, 1145, 1374, 1603, 1832, 2061, 2290, 2519, 2748, 2977, 3206, 3435, 3664, 3893, 4122, 4351, 4580, 4809, 5038, 5267, 5496, 5725, 5954, 6183, 6412, 6641, 6870, 7099, 7328, 7557, 7786, 8015, 8244, 8473, 8702, 8931, 9160, 9389, 9618, 9847, 10076, 10305, 10534, 10763, 10992, 11221, 11450, 11679, 11908, 12137, 12366, 12595, 12824, 13053, 13282, 13511, 13740, 13969, 14198, 14427, 14656, 14885, 15114, 15343, 15572, 15801, 16030, 16259, 16488, 16717, 16946, 17175, 17404, 17633, 17862, 18091, 18320, 18549, 18778, 19007, 19236, 19465, 19694, 19923, 20152, 20381, 20610, 20839, 21068, 21297, 21526, 21755, 21984, 22213, 22442, 22671, 22900, 23129, 23358, 23587, 23816, 24045, 24274, 24503, 24732, 24961, 25190, 25419, 25648, 25877, 26106, 26335, 26564, 26793, 27022, 27251, 27480, 27709, 27938, 28167, 28396, 28625, 28854, 29083, 29312, 29541, 29770, 29999, 30228, 30457, 30686, 30915, 31144, 31373, 31602, 31831, 32060, 32289, 32518, 32747, 32976, 33205, 33434, 33663, 33892, 34121, 34350, 34579, 34808, 35037, 35266, 35495, 35724, 35953, 36182, 36411, 36640, 36869, 37098, 37327, 37556, 37785, 38014, 38243, 38472, 38701, 38930, 39159, 39388, 39617, 39846, 40075, 40304, 40533, 40762, 40991, 41220, 41449, 41678, 41907, 42136, 42365, 42594, 42823, 43052, 43281, 43510, 43739, 43968, 44197, 44426, 44655, 44884, 45113, 45342, 45571, 45800, 46029, 46258, 46487, 46716, 46945, 47174, 47403, 47632, 47861, 48090, 48319, 48548, 48777, 49006, 49235, 49464, 49693, 49922, 50151, 50380, 50609, 50838, 51067, 51296, 51525, 51754, 51983, 52212, 52441, 52670, 52899, 53128, 53357, 53586, 53815, 54044, 54273, 54502, 54731, 54960, 55189, 55418, 55647, 55876, 56105, 56334, 56563, 56792, 57021, 57250, 57479, 57708, 57937, 58166, 58395, 
0, 230, 460, 690, 920, 1150, 1380, 1610, 1840, 2070, 2300, 2530, 2760, 2990, 3220, 3450, 3680, 3910, 4140, 4370, 4600, 4830, 5060, 5290, 5520, 5750, 5980, 6210, 6440, 6670, 6900, 7130, 7360, 7590, 7820, 8050, 8280, 8510, 8740, 8970, 9200, 9430, 9660, 9890, 10120, 10350, 10580, 10810, 11040, 11270, 11500, 11730, 11960, 12190, 12420, 12650, 12880, 13110, 13340, 13570, 13800, 14030, 14260, 14490, 14720, 14950, 15180, 15410, 15640, 15870, 16100, 16330, 16560, 16790, 17020, 17250, 17480, 17710, 17940, 18170, 18400, 18630, 18860, 19090, 19320, 19550, 19780, 20010, 20240, 20470, 20700, 20930, 21160, 21390, 21620, 21850, 22080, 22310, 22540, 22770, 23000, 23230, 23460, 23690, 23920, 24150, 24380, 24610, 24840, 25070, 25300, 25530, 25760, 25990, 26220, 26450, 26680, 26910, 27140, 27370, 27600, 27830, 28060, 28290, 28520, 28750, 28980, 29210, 29440, 29670, 29900, 30130, 30360, 30590, 30820, 31050, 31280, 31510, 31740, 31970, 32200, 32430, 32660, 32890, 33120, 33350, 33580, 33810, 34040, 34270, 34500, 34730, 34960, 35190, 35420, 35650, 35880, 36110, 36340, 36570, 36800, 37030, 37260, 37490, 37720, 37950, 38180, 38410, 38640, 38870, 39100, 39330, 39560, 39790, 40020, 40250, 40480, 40710, 40940, 41170, 41400, 41630, 41860, 42090, 42320, 42550, 42780, 43010, 43240, 43470, 43700, 43930, 44160, 44390, 44620, 44850, 45080, 45310, 45540, 45770, 46000, 46230, 46460, 46690, 46920, 47150, 47380, 47610, 47840, 48070, 48300, 48530, 48760, 48990, 49220, 49450, 49680, 49910, 50140, 50370, 50600, 50830, 51060, 51290, 51520, 51750, 51980, 52210, 52440, 52670, 52900, 53130, 53360, 53590, 53820, 54050, 54280, 54510, 54740, 54970, 55200, 55430, 55660, 55890, 56120, 56350, 56580, 56810, 57040, 57270, 57500, 57730, 57960, 58190, 58420, 58650, 
0, 231, 462, 693, 924, 1155, 1386, 1617, 1848, 2079, 2310, 2541, 2772, 3003, 3234, 3465, 3696, 3927, 4158, 4389, 4620, 4851, 5082, 5313, 5544, 5775, 6006, 6237, 6468, 6699, 6930, 7161, 7392, 7623, 7854, 8085, 8316, 8547, 8778, 9009, 9240, 9471, 9702, 9933, 10164, 10395, 10626, 10857, 11088, 11319, 11550, 11781, 12012, 12243, 12474, 12705, 12936, 13167, 13398, 13629, 13860, 14091, 14322, 14553, 14784, 15015, 15246, 15477, 15708, 15939, 16170, 16401, 16632, 16863, 17094, 17325, 17556, 17787, 18018, 18249, 18480, 18711, 18942, 19173, 19404, 19635, 19866, 20097, 20328, 20559, 20790, 21021, 21252, 21483, 21714, 21945, 22176, 22407, 22638, 22869, 23100, 23331, 23562, 23793, 24024, 24255, 24486, 24717, 24948, 25179, 25410, 25641, 25872, 26103, 26334, 26565, 26796, 27027, 27258, 27489, 27720, 27951, 28182, 28413, 28644, 28875, 29106, 29337, 29568, 29799, 30030, 30261, 30492, 30723, 30954, 31185, 31416, 31647, 31878, 32109, 32340, 32571, 32802, 33033, 33264, 33495, 33726, 33957, 34188, 34419, 34650, 34881, 35112, 35343, 35574, 35805, 36036, 36267, 36498, 36729, 36960, 37191, 37422, 37653, 37884, 38115, 38346, 38577, 38808, 39039, 39270, 39501, 39732, 39963, 40194, 40425, 40656, 40887, 41118, 41349, 41580, 41811, 42042, 42273, 42504, 42735, 42966, 43197, 43428, 43659, 43890, 44121, 44352, 44583, 44814, 45045, 45276, 45507, 45738, 45969, 46200, 46431, 46662, 46893, 47124, 47355, 47586, 47817, 48048, 48279, 48510, 48741, 48972, 49203, 49434, 49665, 49896, 50127, 50358, 50589, 50820, 51051, 51282, 51513, 51744, 51975, 52206, 52437, 52668, 52899, 53130, 53361, 53592, 53823, 54054, 54285, 54516, 54747, 54978, 55209, 55440, 55671, 55902, 56133, 56364, 56595, 56826, 57057, 57288, 57519, 57750, 57981, 58212, 58443, 58674, 58905, 
0, 232, 464, 696, 928, 1160, 1392, 1624, 1856, 2088, 2320, 2552, 2784, 3016, 3248, 3480, 3712, 3944, 4176, 4408, 4640, 4872, 5104, 5336, 5568, 5800, 6032, 6264, 6496, 6728, 6960, 7192, 7424, 7656, 7888, 8120, 8352, 8584, 8816, 9048, 9280, 9512, 9744, 9976, 10208, 10440, 10672, 10904, 11136, 11368, 11600, 11832, 12064, 12296, 12528, 12760, 12992, 13224, 13456, 13688, 13920, 14152, 14384, 14616, 14848, 15080, 15312, 15544, 15776, 16008, 16240, 16472, 16704, 16936, 17168, 17400, 17632, 17864, 18096, 18328, 18560, 18792, 19024, 19256, 19488, 19720, 19952, 20184, 20416, 20648, 20880, 21112, 21344, 21576, 21808, 22040, 22272, 22504, 22736, 22968, 23200, 23432, 23664, 23896, 24128, 24360, 24592, 24824, 25056, 25288, 25520, 25752, 25984, 26216, 26448, 26680, 26912, 27144, 27376, 27608, 27840, 28072, 28304, 28536, 28768, 29000, 29232, 29464, 29696, 29928, 30160, 30392, 30624, 30856, 31088, 31320, 31552, 31784, 32016, 32248, 32480, 32712, 32944, 33176, 33408, 33640, 33872, 34104, 34336, 34568, 34800, 35032, 35264, 35496, 35728, 35960, 36192, 36424, 36656, 36888, 37120, 37352, 37584, 37816, 38048, 38280, 38512, 38744, 38976, 39208, 39440, 39672, 39904, 40136, 40368, 40600, 40832, 41064, 41296, 41528, 41760, 41992, 42224, 42456, 42688, 42920, 43152, 43384, 43616, 43848, 44080, 44312, 44544, 44776, 45008, 45240, 45472, 45704, 45936, 46168, 46400, 46632, 46864, 47096, 47328, 47560, 47792, 48024, 48256, 48488, 48720, 48952, 49184, 49416, 49648, 49880, 50112, 50344, 50576, 50808, 51040, 51272, 51504, 51736, 51968, 52200, 52432, 52664, 52896, 53128, 53360, 53592, 53824, 54056, 54288, 54520, 54752, 54984, 55216, 55448, 55680, 55912, 56144, 56376, 56608, 56840, 57072, 57304, 57536, 57768, 58000, 58232, 58464, 58696, 58928, 59160, 
0, 233, 466, 699, 932, 1165, 1398, 1631, 1864, 2097, 2330, 2563, 2796, 3029, 3262, 3495, 3728, 3961, 4194, 4427, 4660, 4893, 5126, 5359, 5592, 5825, 6058, 6291, 6524, 6757, 6990, 7223, 7456, 7689, 7922, 8155, 8388, 8621, 8854, 9087, 9320, 9553, 9786, 10019, 10252, 10485, 10718, 10951, 11184, 11417, 11650, 11883, 12116, 12349, 12582, 12815, 13048, 13281, 13514, 13747, 13980, 14213, 14446, 14679, 14912, 15145, 15378, 15611, 15844, 16077, 16310, 16543, 16776, 17009, 17242, 17475, 17708, 17941, 18174, 18407, 18640, 18873, 19106, 19339, 19572, 19805, 20038, 20271, 20504, 20737, 20970, 21203, 21436, 21669, 21902, 22135, 22368, 22601, 22834, 23067, 23300, 23533, 23766, 23999, 24232, 24465, 24698, 24931, 25164, 25397, 25630, 25863, 26096, 26329, 26562, 26795, 27028, 27261, 27494, 27727, 27960, 28193, 28426, 28659, 28892, 29125, 29358, 29591, 29824, 30057, 30290, 30523, 30756, 30989, 31222, 31455, 31688, 31921, 32154, 32387, 32620, 32853, 33086, 33319, 33552, 33785, 34018, 34251, 34484, 34717, 34950, 35183, 35416, 35649, 35882, 36115, 36348, 36581, 36814, 37047, 37280, 37513, 37746, 37979, 38212, 38445, 38678, 38911, 39144, 39377, 39610, 39843, 40076, 40309, 40542, 40775, 41008, 41241, 41474, 41707, 41940, 42173, 42406, 42639, 42872, 43105, 43338, 43571, 43804, 44037, 44270, 44503, 44736, 44969, 45202, 45435, 45668, 45901, 46134, 46367, 46600, 46833, 47066, 47299, 47532, 47765, 47998, 48231, 48464, 48697, 48930, 49163, 49396, 49629, 49862, 50095, 50328, 50561, 50794, 51027, 51260, 51493, 51726, 51959, 52192, 52425, 52658, 52891, 53124, 53357, 53590, 53823, 54056, 54289, 54522, 54755, 54988, 55221, 55454, 55687, 55920, 56153, 56386, 56619, 56852, 57085, 57318, 57551, 57784, 58017, 58250, 58483, 58716, 58949, 59182, 59415, 
0, 234, 468, 702, 936, 1170, 1404, 1638, 1872, 2106, 2340, 2574, 2808, 3042, 3276, 3510, 3744, 3978, 4212, 4446, 4680, 4914, 5148, 5382, 5616, 5850, 6084, 6318, 6552, 6786, 7020, 7254, 7488, 7722, 7956, 8190, 8424, 8658, 8892, 9126, 9360, 9594, 9828, 10062, 10296, 10530, 10764, 10998, 11232, 11466, 11700, 11934, 12168, 12402, 12636, 12870, 13104, 13338, 13572, 13806, 14040, 14274, 14508, 14742, 14976, 15210, 15444, 15678, 15912, 16146, 16380, 16614, 16848, 17082, 17316, 17550, 17784, 18018, 18252, 18486, 18720, 18954, 19188, 19422, 19656, 19890, 20124, 20358, 20592, 20826, 21060, 21294, 21528, 21762, 21996, 22230, 22464, 22698, 22932, 23166, 23400, 23634, 23868, 24102, 24336, 24570, 24804, 25038, 25272, 25506, 25740, 25974, 26208, 26442, 26676, 26910, 27144, 27378, 27612, 27846, 28080, 28314, 28548, 28782, 29016, 29250, 29484, 29718, 29952, 30186, 30420, 30654, 30888, 31122, 31356, 31590, 31824, 32058, 32292, 32526, 32760, 32994, 33228, 33462, 33696, 33930, 34164, 34398, 34632, 34866, 35100, 35334, 35568, 35802, 36036, 36270, 36504, 36738, 36972, 37206, 37440, 37674, 37908, 38142, 38376, 38610, 38844, 39078, 39312, 39546, 39780, 40014, 40248, 40482, 40716, 40950, 41184, 41418, 41652, 41886, 42120, 42354, 42588, 42822, 43056, 43290, 43524, 43758, 43992, 44226, 44460, 44694, 44928, 45162, 45396, 45630, 45864, 46098, 46332, 46566, 46800, 47034, 47268, 47502, 47736, 47970, 48204, 48438, 48672, 48906, 49140, 49374, 49608, 49842, 50076, 50310, 50544, 50778, 51012, 51246, 51480, 51714, 51948, 52182, 52416, 52650, 52884, 53118, 53352, 53586, 53820, 54054, 54288, 54522, 54756, 54990, 55224, 55458, 55692, 55926, 56160, 56394, 56628, 56862, 57096, 57330, 57564, 57798, 58032, 58266, 58500, 58734, 58968, 59202, 59436, 59670, 
0, 235, 470, 705, 940, 1175, 1410, 1645, 1880, 2115, 2350, 2585, 2820, 3055, 3290, 3525, 3760, 3995, 4230, 4465, 4700, 4935, 5170, 5405, 5640, 5875, 6110, 6345, 6580, 6815, 7050, 7285, 7520, 7755, 7990, 8225, 8460, 8695, 8930, 9165, 9400, 9635, 9870, 10105, 10340, 10575, 10810, 11045, 11280, 11515, 11750, 11985, 12220, 12455, 12690, 12925, 13160, 13395, 13630, 13865, 14100, 14335, 14570, 14805, 15040, 15275, 15510, 15745, 15980, 16215, 16450, 16685, 16920, 17155, 17390, 17625, 17860, 18095, 18330, 18565, 18800, 19035, 19270, 19505, 19740, 19975, 20210, 20445, 20680, 20915, 21150, 21385, 21620, 21855, 22090, 22325, 22560, 22795, 23030, 23265, 23500, 23735, 23970, 24205, 24440, 24675, 24910, 25145, 25380, 25615, 25850, 26085, 26320, 26555, 26790, 27025, 27260, 27495, 27730, 27965, 28200, 28435, 28670, 28905, 29140, 29375, 29610, 29845, 30080, 30315, 30550, 30785, 31020, 31255, 31490, 31725, 31960, 32195, 32430, 32665, 32900, 33135, 33370, 33605, 33840, 34075, 34310, 34545, 34780, 35015, 35250, 35485, 35720, 35955, 36190, 36425, 36660, 36895, 37130, 37365, 37600, 37835, 38070, 38305, 38540, 38775, 39010, 39245, 39480, 39715, 39950, 40185, 40420, 40655, 40890, 41125, 41360, 41595, 41830, 42065, 42300, 42535, 42770, 43005, 43240, 43475, 43710, 43945, 44180, 44415, 44650, 44885, 45120, 45355, 45590, 45825, 46060, 46295, 46530, 46765, 47000, 47235, 47470, 47705, 47940, 48175, 48410, 48645, 48880, 49115, 49350, 49585, 49820, 50055, 50290, 50525, 50760, 50995, 51230, 51465, 51700, 51935, 52170, 52405, 52640, 52875, 53110, 53345, 53580, 53815, 54050, 54285, 54520, 54755, 54990, 55225, 55460, 55695, 55930, 56165, 56400, 56635, 56870, 57105, 57340, 57575, 57810, 58045, 58280, 58515, 58750, 58985, 59220, 59455, 59690, 59925, 
0, 236, 472, 708, 944, 1180, 1416, 1652, 1888, 2124, 2360, 2596, 2832, 3068, 3304, 3540, 3776, 4012, 4248, 4484, 4720, 4956, 5192, 5428, 5664, 5900, 6136, 6372, 6608, 6844, 7080, 7316, 7552, 7788, 8024, 8260, 8496, 8732, 8968, 9204, 9440, 9676, 9912, 10148, 10384, 10620, 10856, 11092, 11328, 11564, 11800, 12036, 12272, 12508, 12744, 12980, 13216, 13452, 13688, 13924, 14160, 14396, 14632, 14868, 15104, 15340, 15576, 15812, 16048, 16284, 16520, 16756, 16992, 17228, 17464, 17700, 17936, 18172, 18408, 18644, 18880, 19116, 19352, 19588, 19824, 20060, 20296, 20532, 20768, 21004, 21240, 21476, 21712, 21948, 22184, 22420, 22656, 22892, 23128, 23364, 23600, 23836, 24072, 24308, 24544, 24780, 25016, 25252, 25488, 25724, 25960, 26196, 26432, 26668, 26904, 27140, 27376, 27612, 27848, 28084, 28320, 28556, 28792, 29028, 29264, 29500, 29736, 29972, 30208, 30444, 30680, 30916, 31152, 31388, 31624, 31860, 32096, 32332, 32568, 32804, 33040, 33276, 33512, 33748, 33984, 34220, 34456, 34692, 34928, 35164, 35400, 35636, 35872, 36108, 36344, 36580, 36816, 37052, 37288, 37524, 37760, 37996, 38232, 38468, 38704, 38940, 39176, 39412, 39648, 39884, 40120, 40356, 40592, 40828, 41064, 41300, 41536, 41772, 42008, 42244, 42480, 42716, 42952, 43188, 43424, 43660, 43896, 44132, 44368, 44604, 44840, 45076, 45312, 45548, 45784, 46020, 46256, 46492, 46728, 46964, 47200, 47436, 47672, 47908, 48144, 48380, 48616, 48852, 49088, 49324, 49560, 49796, 50032, 50268, 50504, 50740, 50976, 51212, 51448, 51684, 51920, 52156, 52392, 52628, 52864, 53100, 53336, 53572, 53808, 54044, 54280, 54516, 54752, 54988, 55224, 55460, 55696, 55932, 56168, 56404, 56640, 56876, 57112, 57348, 57584, 57820, 58056, 58292, 58528, 58764, 59000, 59236, 59472, 59708, 59944, 60180, 
0, 237, 474, 711, 948, 1185, 1422, 1659, 1896, 2133, 2370, 2607, 2844, 3081, 3318, 3555, 3792, 4029, 4266, 4503, 4740, 4977, 5214, 5451, 5688, 5925, 6162, 6399, 6636, 6873, 7110, 7347, 7584, 7821, 8058, 8295, 8532, 8769, 9006, 9243, 9480, 9717, 9954, 10191, 10428, 10665, 10902, 11139, 11376, 11613, 11850, 12087, 12324, 12561, 12798, 13035, 13272, 13509, 13746, 13983, 14220, 14457, 14694, 14931, 15168, 15405, 15642, 15879, 16116, 16353, 16590, 16827, 17064, 17301, 17538, 17775, 18012, 18249, 18486, 18723, 18960, 19197, 19434, 19671, 19908, 20145, 20382, 20619, 20856, 21093, 21330, 21567, 21804, 22041, 22278, 22515, 22752, 22989, 23226, 23463, 23700, 23937, 24174, 24411, 24648, 24885, 25122, 25359, 25596, 25833, 26070, 26307, 26544, 26781, 27018, 27255, 27492, 27729, 27966, 28203, 28440, 28677, 28914, 29151, 29388, 29625, 29862, 30099, 30336, 30573, 30810, 31047, 31284, 31521, 31758, 31995, 32232, 32469, 32706, 32943, 33180, 33417, 33654, 33891, 34128, 34365, 34602, 34839, 35076, 35313, 35550, 35787, 36024, 36261, 36498, 36735, 36972, 37209, 37446, 37683, 37920, 38157, 38394, 38631, 38868, 39105, 39342, 39579, 39816, 40053, 40290, 40527, 40764, 41001, 41238, 41475, 41712, 41949, 42186, 42423, 42660, 42897, 43134, 43371, 43608, 43845, 44082, 44319, 44556, 44793, 45030, 45267, 45504, 45741, 45978, 46215, 46452, 46689, 46926, 47163, 47400, 47637, 47874, 48111, 48348, 48585, 48822, 49059, 49296, 49533, 49770, 50007, 50244, 50481, 50718, 50955, 51192, 51429, 51666, 51903, 52140, 52377, 52614, 52851, 53088, 53325, 53562, 53799, 54036, 54273, 54510, 54747, 54984, 55221, 55458, 55695, 55932, 56169, 56406, 56643, 56880, 57117, 57354, 57591, 57828, 58065, 58302, 58539, 58776, 59013, 59250, 59487, 59724, 59961, 60198, 60435, 
0, 238, 476, 714, 952, 1190, 1428, 1666, 1904, 2142, 2380, 2618, 2856, 3094, 3332, 3570, 3808, 4046, 4284, 4522, 4760, 4998, 5236, 5474, 5712, 5950, 6188, 6426, 6664, 6902, 7140, 7378, 7616, 7854, 8092, 8330, 8568, 8806, 9044, 9282, 9520, 9758, 9996, 10234, 10472, 10710, 10948, 11186, 11424, 11662, 11900, 12138, 12376, 12614, 12852, 13090, 13328, 13566, 13804, 14042, 14280, 14518, 14756, 14994, 15232, 15470, 15708, 15946, 16184, 16422, 16660, 16898, 17136, 17374, 17612, 17850, 18088, 18326, 18564, 18802, 19040, 19278, 19516, 19754, 19992, 20230, 20468, 20706, 20944, 21182, 21420, 21658, 21896, 22134, 22372, 22610, 22848, 23086, 23324, 23562, 23800, 24038, 24276, 24514, 24752, 24990, 25228, 25466, 25704, 25942, 26180, 26418, 26656, 26894, 27132, 27370, 27608, 27846, 28084, 28322, 28560, 28798, 29036, 29274, 29512, 29750, 29988, 30226, 30464, 30702, 30940, 31178, 31416, 31654, 31892, 32130, 32368, 32606, 32844, 33082, 33320, 33558, 33796, 34034, 34272, 34510, 34748, 34986, 35224, 35462, 35700, 35938, 36176, 36414, 36652, 36890, 37128, 37366, 37604, 37842, 38080, 38318, 38556, 38794, 39032, 39270, 39508, 39746, 39984, 40222, 40460, 40698, 40936, 41174, 41412, 41650, 41888, 42126, 42364, 42602, 42840, 43078, 43316, 43554, 43792, 44030, 44268, 44506, 44744, 44982, 45220, 45458, 45696, 45934, 46172, 46410, 46648, 46886, 47124, 47362, 47600, 47838, 48076, 48314, 48552, 48790, 49028, 49266, 49504, 49742, 49980, 50218, 50456, 50694, 50932, 51170, 51408, 51646, 51884, 52122, 52360, 52598, 52836, 53074, 53312, 53550, 53788, 54026, 54264, 54502, 54740, 54978, 55216, 55454, 55692, 55930, 56168, 56406, 56644, 56882, 57120, 57358, 57596, 57834, 58072, 58310, 58548, 58786, 59024, 59262, 59500, 59738, 59976, 60214, 60452, 60690, 
0, 239, 478, 717, 956, 1195, 1434, 1673, 1912, 2151, 2390, 2629, 2868, 3107, 3346, 3585, 3824, 4063, 4302, 4541, 4780, 5019, 5258, 5497, 5736, 5975, 6214, 6453, 6692, 6931, 7170, 7409, 7648, 7887, 8126, 8365, 8604, 8843, 9082, 9321, 9560, 9799, 10038, 10277, 10516, 10755, 10994, 11233, 11472, 11711, 11950, 12189, 12428, 12667, 12906, 13145, 13384, 13623, 13862, 14101, 14340, 14579, 14818, 15057, 15296, 15535, 15774, 16013, 16252, 16491, 16730, 16969, 17208, 17447, 17686, 17925, 18164, 18403, 18642, 18881, 19120, 19359, 19598, 19837, 20076, 20315, 20554, 20793, 21032, 21271, 21510, 21749, 21988, 22227, 22466, 22705, 22944, 23183, 23422, 23661, 23900, 24139, 24378, 24617, 24856, 25095, 25334, 25573, 25812, 26051, 26290, 26529, 26768, 27007, 27246, 27485, 27724, 27963, 28202, 28441, 28680, 28919, 29158, 29397, 29636, 29875, 30114, 30353, 30592, 30831, 31070, 31309, 31548, 31787, 32026, 32265, 32504, 32743, 32982, 33221, 33460, 33699, 33938, 34177, 34416, 34655, 34894, 35133, 35372, 35611, 35850, 36089, 36328, 36567, 36806, 37045, 37284, 37523, 37762, 38001, 38240, 38479, 38718, 38957, 39196, 39435, 39674, 39913, 40152, 40391, 40630, 40869, 41108, 41347, 41586, 41825, 42064, 42303, 42542, 42781, 43020, 43259, 43498, 43737, 43976, 44215, 44454, 44693, 44932, 45171, 45410, 45649, 45888, 46127, 46366, 46605, 46844, 47083, 47322, 47561, 47800, 48039, 48278, 48517, 48756, 48995, 49234, 49473, 49712, 49951, 50190, 50429, 50668, 50907, 51146, 51385, 51624, 51863, 52102, 52341, 52580, 52819, 53058, 53297, 53536, 53775, 54014, 54253, 54492, 54731, 54970, 55209, 55448, 55687, 55926, 56165, 56404, 56643, 56882, 57121, 57360, 57599, 57838, 58077, 58316, 58555, 58794, 59033, 59272, 59511, 59750, 59989, 60228, 60467, 60706, 60945, 
0, 240, 480, 720, 960, 1200, 1440, 1680, 1920, 2160, 2400, 2640, 2880, 3120, 3360, 3600, 3840, 4080, 4320, 4560, 4800, 5040, 5280, 5520, 5760, 6000, 6240, 6480, 6720, 6960, 7200, 7440, 7680, 7920, 8160, 8400, 8640, 8880, 9120, 9360, 9600, 9840, 10080, 10320, 10560, 10800, 11040, 11280, 11520, 11760, 12000, 12240, 12480, 12720, 12960, 13200, 13440, 13680, 13920, 14160, 14400, 14640, 14880, 15120, 15360, 15600, 15840, 16080, 16320, 16560, 16800, 17040, 17280, 17520, 17760, 18000, 18240, 18480, 18720, 18960, 19200, 19440, 19680, 19920, 20160, 20400, 20640, 20880, 21120, 21360, 21600, 21840, 22080, 22320, 22560, 22800, 23040, 23280, 23520, 23760, 24000, 24240, 24480, 24720, 24960, 25200, 25440, 25680, 25920, 26160, 26400, 26640, 26880, 27120, 27360, 27600, 27840, 28080, 28320, 28560, 28800, 29040, 29280, 29520, 29760, 30000, 30240, 30480, 30720, 30960, 31200, 31440, 31680, 31920, 32160, 32400, 32640, 32880, 33120, 33360, 33600, 33840, 34080, 34320, 34560, 34800, 35040, 35280, 35520, 35760, 36000, 36240, 36480, 36720, 36960, 37200, 37440, 37680, 37920, 38160, 38400, 38640, 38880, 39120, 39360, 39600, 39840, 40080, 40320, 40560, 40800, 41040, 41280, 41520, 41760, 42000, 42240, 42480, 42720, 42960, 43200, 43440, 43680, 43920, 44160, 44400, 44640, 44880, 45120, 45360, 45600, 45840, 46080, 46320, 46560, 46800, 47040, 47280, 47520, 47760, 48000, 48240, 48480, 48720, 48960, 49200, 49440, 49680, 49920, 50160, 50400, 50640, 50880, 51120, 51360, 51600, 51840, 52080, 52320, 52560, 52800, 53040, 53280, 53520, 53760, 54000, 54240, 54480, 54720, 54960, 55200, 55440, 55680, 55920, 56160, 56400, 56640, 56880, 57120, 57360, 57600, 57840, 58080, 58320, 58560, 58800, 59040, 59280, 59520, 59760, 60000, 60240, 60480, 60720, 60960, 61200, 
0, 241, 482, 723, 964, 1205, 1446, 1687, 1928, 2169, 2410, 2651, 2892, 3133, 3374, 3615, 3856, 4097, 4338, 4579, 4820, 5061, 5302, 5543, 5784, 6025, 6266, 6507, 6748, 6989, 7230, 7471, 7712, 7953, 8194, 8435, 8676, 8917, 9158, 9399, 9640, 9881, 10122, 10363, 10604, 10845, 11086, 11327, 11568, 11809, 12050, 12291, 12532, 12773, 13014, 13255, 13496, 13737, 13978, 14219, 14460, 14701, 14942, 15183, 15424, 15665, 15906, 16147, 16388, 16629, 16870, 17111, 17352, 17593, 17834, 18075, 18316, 18557, 18798, 19039, 19280, 19521, 19762, 20003, 20244, 20485, 20726, 20967, 21208, 21449, 21690, 21931, 22172, 22413, 22654, 22895, 23136, 23377, 23618, 23859, 24100, 24341, 24582, 24823, 25064, 25305, 25546, 25787, 26028, 26269, 26510, 26751, 26992, 27233, 27474, 27715, 27956, 28197, 28438, 28679, 28920, 29161, 29402, 29643, 29884, 30125, 30366, 30607, 30848, 31089, 31330, 31571, 31812, 32053, 32294, 32535, 32776, 33017, 33258, 33499, 33740, 33981, 34222, 34463, 34704, 34945, 35186, 35427, 35668, 35909, 36150, 36391, 36632, 36873, 37114, 37355, 37596, 37837, 38078, 38319, 38560, 38801, 39042, 39283, 39524, 39765, 40006, 40247, 40488, 40729, 40970, 41211, 41452, 41693, 41934, 42175, 42416, 42657, 42898, 43139, 43380, 43621, 43862, 44103, 44344, 44585, 44826, 45067, 45308, 45549, 45790, 46031, 46272, 46513, 46754, 46995, 47236, 47477, 47718, 47959, 48200, 48441, 48682, 48923, 49164, 49405, 49646, 49887, 50128, 50369, 50610, 50851, 51092, 51333, 51574, 51815, 52056, 52297, 52538, 52779, 53020, 53261, 53502, 53743, 53984, 54225, 54466, 54707, 54948, 55189, 55430, 55671, 55912, 56153, 56394, 56635, 56876, 57117, 57358, 57599, 57840, 58081, 58322, 58563, 58804, 59045, 59286, 59527, 59768, 60009, 60250, 60491, 60732, 60973, 61214, 61455, 
0, 242, 484, 726, 968, 1210, 1452, 1694, 1936, 2178, 2420, 2662, 2904, 3146, 3388, 3630, 3872, 4114, 4356, 4598, 4840, 5082, 5324, 5566, 5808, 6050, 6292, 6534, 6776, 7018, 7260, 7502, 7744, 7986, 8228, 8470, 8712, 8954, 9196, 9438, 9680, 9922, 10164, 10406, 10648, 10890, 11132, 11374, 11616, 11858, 12100, 12342, 12584, 12826, 13068, 13310, 13552, 13794, 14036, 14278, 14520, 14762, 15004, 15246, 15488, 15730, 15972, 16214, 16456, 16698, 16940, 17182, 17424, 17666, 17908, 18150, 18392, 18634, 18876, 19118, 19360, 19602, 19844, 20086, 20328, 20570, 20812, 21054, 21296, 21538, 21780, 22022, 22264, 22506, 22748, 22990, 23232, 23474, 23716, 23958, 24200, 24442, 24684, 24926, 25168, 25410, 25652, 25894, 26136, 26378, 26620, 26862, 27104, 27346, 27588, 27830, 28072, 28314, 28556, 28798, 29040, 29282, 29524, 29766, 30008, 30250, 30492, 30734, 30976, 31218, 31460, 31702, 31944, 32186, 32428, 32670, 32912, 33154, 33396, 33638, 33880, 34122, 34364, 34606, 34848, 35090, 35332, 35574, 35816, 36058, 36300, 36542, 36784, 37026, 37268, 37510, 37752, 37994, 38236, 38478, 38720, 38962, 39204, 39446, 39688, 39930, 40172, 40414, 40656, 40898, 41140, 41382, 41624, 41866, 42108, 42350, 42592, 42834, 43076, 43318, 43560, 43802, 44044, 44286, 44528, 44770, 45012, 45254, 45496, 45738, 45980, 46222, 46464, 46706, 46948, 47190, 47432, 47674, 47916, 48158, 48400, 48642, 48884, 49126, 49368, 49610, 49852, 50094, 50336, 50578, 50820, 51062, 51304, 51546, 51788, 52030, 52272, 52514, 52756, 52998, 53240, 53482, 53724, 53966, 54208, 54450, 54692, 54934, 55176, 55418, 55660, 55902, 56144, 56386, 56628, 56870, 57112, 57354, 57596, 57838, 58080, 58322, 58564, 58806, 59048, 59290, 59532, 59774, 60016, 60258, 60500, 60742, 60984, 61226, 61468, 61710, 
0, 243, 486, 729, 972, 1215, 1458, 1701, 1944, 2187, 2430, 2673, 2916, 3159, 3402, 3645, 3888, 4131, 4374, 4617, 4860, 5103, 5346, 5589, 5832, 6075, 6318, 6561, 6804, 7047, 7290, 7533, 7776, 8019, 8262, 8505, 8748, 8991, 9234, 9477, 9720, 9963, 10206, 10449, 10692, 10935, 11178, 11421, 11664, 11907, 12150, 12393, 12636, 12879, 13122, 13365, 13608, 13851, 14094, 14337, 14580, 14823, 15066, 15309, 15552, 15795, 16038, 16281, 16524, 16767, 17010, 17253, 17496, 17739, 17982, 18225, 18468, 18711, 18954, 19197, 19440, 19683, 19926, 20169, 20412, 20655, 20898, 21141, 21384, 21627, 21870, 22113, 22356, 22599, 22842, 23085, 23328, 23571, 23814, 24057, 24300, 24543, 24786, 25029, 25272, 25515, 25758, 26001, 26244, 26487, 26730, 26973, 27216, 27459, 27702, 27945, 28188, 28431, 28674, 28917, 29160, 29403, 29646, 29889, 30132, 30375, 30618, 30861, 31104, 31347, 31590, 31833, 32076, 32319, 32562, 32805, 33048, 33291, 33534, 33777, 34020, 34263, 34506, 34749, 34992, 35235, 35478, 35721, 35964, 36207, 36450, 36693, 36936, 37179, 37422, 37665, 37908, 38151, 38394, 38637, 38880, 39123, 39366, 39609, 39852, 40095, 40338, 40581, 40824, 41067, 41310, 41553, 41796, 42039, 42282, 42525, 42768, 43011, 43254, 43497, 43740, 43983, 44226, 44469, 44712, 44955, 45198, 45441, 45684, 45927, 46170, 46413, 46656, 46899, 47142, 47385, 47628, 47871, 48114, 48357, 48600, 48843, 49086, 49329, 49572, 49815, 50058, 50301, 50544, 50787, 51030, 51273, 51516, 51759, 52002, 52245, 52488, 52731, 52974, 53217, 53460, 53703, 53946, 54189, 54432, 54675, 54918, 55161, 55404, 55647, 55890, 56133, 56376, 56619, 56862, 57105, 57348, 57591, 57834, 58077, 58320, 58563, 58806, 59049, 59292, 59535, 59778, 60021, 60264, 60507, 60750, 60993, 61236, 61479, 61722, 61965, 
0, 244, 488, 732, 976, 1220, 1464, 1708, 1952, 2196, 2440, 2684, 2928, 3172, 3416, 3660, 3904, 4148, 4392, 4636, 4880, 5124, 5368, 5612, 5856, 6100, 6344, 6588, 6832, 7076, 7320, 7564, 7808, 8052, 8296, 8540, 8784, 9028, 9272, 9516, 9760, 10004, 10248, 10492, 10736, 10980, 11224, 11468, 11712, 11956, 12200, 12444, 12688, 12932, 13176, 13420, 13664, 13908, 14152, 14396, 14640, 14884, 15128, 15372, 15616, 15860, 16104, 16348, 16592, 16836, 17080, 17324, 17568, 17812, 18056, 18300, 18544, 18788, 19032, 19276, 19520, 19764, 20008, 20252, 20496, 20740, 20984, 21228, 21472, 21716, 21960, 22204, 22448, 22692, 22936, 23180, 23424, 23668, 23912, 24156, 24400, 24644, 24888, 25132, 25376, 25620, 25864, 26108, 26352, 26596, 26840, 27084, 27328, 27572, 27816, 28060, 28304, 28548, 28792, 29036, 29280, 29524, 29768, 30012, 30256, 30500, 30744, 30988, 31232, 31476, 31720, 31964, 32208, 32452, 32696, 32940, 33184, 33428, 33672, 33916, 34160, 34404, 34648, 34892, 35136, 35380, 35624, 35868, 36112, 36356, 36600, 36844, 37088, 37332, 37576, 37820, 38064, 38308, 38552, 38796, 39040, 39284, 39528, 39772, 40016, 40260, 40504, 40748, 40992, 41236, 41480, 41724, 41968, 42212, 42456, 42700, 42944, 43188, 43432, 43676, 43920, 44164, 44408, 44652, 44896, 45140, 45384, 45628, 45872, 46116, 46360, 46604, 46848, 47092, 47336, 47580, 47824, 48068, 48312, 48556, 48800, 49044, 49288, 49532, 49776, 50020, 50264, 50508, 50752, 50996, 51240, 51484, 51728, 51972, 52216, 52460, 52704, 52948, 53192, 53436, 53680, 53924, 54168, 54412, 54656, 54900, 55144, 55388, 55632, 55876, 56120, 56364, 56608, 56852, 57096, 57340, 57584, 57828, 58072, 58316, 58560, 58804, 59048, 59292, 59536, 59780, 60024, 60268, 60512, 60756, 61000, 61244, 61488, 61732, 61976, 62220, 
0, 245, 490, 735, 980, 1225, 1470, 1715, 1960, 2205, 2450, 2695, 2940, 3185, 3430, 3675, 3920, 4165, 4410, 4655, 4900, 5145, 5390, 5635, 5880, 6125, 6370, 6615, 6860, 7105, 7350, 7595, 7840, 8085, 8330, 8575, 8820, 9065, 9310, 9555, 9800, 10045, 10290, 10535, 10780, 11025, 11270, 11515, 11760, 12005, 12250, 12495, 12740, 12985, 13230, 13475, 13720, 13965, 14210, 14455, 14700, 14945, 15190, 15435, 15680, 15925, 16170, 16415, 16660, 16905, 17150, 17395, 17640, 17885, 18130, 18375, 18620, 18865, 19110, 19355, 19600, 19845, 20090, 20335, 20580, 20825, 21070, 21315, 21560, 21805, 22050, 22295, 22540, 22785, 23030, 23275, 23520, 23765, 24010, 24255, 24500, 24745, 24990, 25235, 25480, 25725, 25970, 26215, 26460, 26705, 26950, 27195, 27440, 27685, 27930, 28175, 28420, 28665, 28910, 29155, 29400, 29645, 29890, 30135, 30380, 30625, 30870, 31115, 31360, 31605, 31850, 32095, 32340, 32585, 32830, 33075, 33320, 33565, 33810, 34055, 34300, 34545, 34790, 35035, 35280, 35525, 35770, 36015, 36260, 36505, 36750, 36995, 37240, 37485, 37730, 37975, 38220, 38465, 38710, 38955, 39200, 39445, 39690, 39935, 40180, 40425, 40670, 40915, 41160, 41405, 41650, 41895, 42140, 42385, 42630, 42875, 43120, 43365, 43610, 43855, 44100, 44345, 44590, 44835, 45080, 45325, 45570, 45815, 46060, 46305, 46550, 46795, 47040, 47285, 47530, 47775, 48020, 48265, 48510, 48755, 49000, 49245, 49490, 49735, 49980, 50225, 50470, 50715, 50960, 51205, 51450, 51695, 51940, 52185, 52430, 52675, 52920, 53165, 53410, 53655, 53900, 54145, 54390, 54635, 54880, 55125, 55370, 55615, 55860, 56105, 56350, 56595, 56840, 57085, 57330, 57575, 57820, 58065, 58310, 58555, 58800, 59045, 59290, 59535, 59780, 60025, 60270, 60515, 60760, 61005, 61250, 61495, 61740, 61985, 62230, 62475, 
0, 246, 492, 738, 984, 1230, 1476, 1722, 1968, 2214, 2460, 2706, 2952, 3198, 3444, 3690, 3936, 4182, 4428, 4674, 4920, 5166, 5412, 5658, 5904, 6150, 6396, 6642, 6888, 7134, 7380, 7626, 7872, 8118, 8364, 8610, 8856, 9102, 9348, 9594, 9840, 10086, 10332, 10578, 10824, 11070, 11316, 11562, 11808, 12054, 12300, 12546, 12792, 13038, 13284, 13530, 13776, 14022, 14268, 14514, 14760, 15006, 15252, 15498, 15744, 15990, 16236, 16482, 16728, 16974, 17220, 17466, 17712, 17958, 18204, 18450, 18696, 18942, 19188, 19434, 19680, 19926, 20172, 20418, 20664, 20910, 21156, 21402, 21648, 21894, 22140, 22386, 22632, 22878, 23124, 23370, 23616, 23862, 24108, 24354, 24600, 24846, 25092, 25338, 25584, 25830, 26076, 26322, 26568, 26814, 27060, 27306, 27552, 27798, 28044, 28290, 28536, 28782, 29028, 29274, 29520, 29766, 30012, 30258, 30504, 30750, 30996, 31242, 31488, 31734, 31980, 32226, 32472, 32718, 32964, 33210, 33456, 33702, 33948, 34194, 34440, 34686, 34932, 35178, 35424, 35670, 35916, 36162, 36408, 36654, 36900, 37146, 37392, 37638, 37884, 38130, 38376, 38622, 38868, 39114, 39360, 39606, 39852, 40098, 40344, 40590, 40836, 41082, 41328, 41574, 41820, 42066, 42312, 42558, 42804, 43050, 43296, 43542, 43788, 44034, 44280, 44526, 44772, 45018, 45264, 45510, 45756, 46002, 46248, 46494, 46740, 46986, 47232, 47478, 47724, 47970, 48216, 48462, 48708, 48954, 49200, 49446, 49692, 49938, 50184, 50430, 50676, 50922, 51168, 51414, 51660, 51906, 52152, 52398, 52644, 52890, 53136, 53382, 53628, 53874, 54120, 54366, 54612, 54858, 55104, 55350, 55596, 55842, 56088, 56334, 56580, 56826, 57072, 57318, 57564, 57810, 58056, 58302, 58548, 58794, 59040, 59286, 59532, 59778, 60024, 60270, 60516, 60762, 61008, 61254, 61500, 61746, 61992, 62238, 62484, 62730, 
0, 247, 494, 741, 988, 1235, 1482, 1729, 1976, 2223, 2470, 2717, 2964, 3211, 3458, 3705, 3952, 4199, 4446, 4693, 4940, 5187, 5434, 5681, 5928, 6175, 6422, 6669, 6916, 7163, 7410, 7657, 7904, 8151, 8398, 8645, 8892, 9139, 9386, 9633, 9880, 10127, 10374, 10621, 10868, 11115, 11362, 11609, 11856, 12103, 12350, 12597, 12844, 13091, 13338, 13585, 13832, 14079, 14326, 14573, 14820, 15067, 15314, 15561, 15808, 16055, 16302, 16549, 16796, 17043, 17290, 17537, 17784, 18031, 18278, 18525, 18772, 19019, 19266, 19513, 19760, 20007, 20254, 20501, 20748, 20995, 21242, 21489, 21736, 21983, 22230, 22477, 22724, 22971, 23218, 23465, 23712, 23959, 24206, 24453, 24700, 24947, 25194, 25441, 25688, 25935, 26182, 26429, 26676, 26923, 27170, 27417, 27664, 27911, 28158, 28405, 28652, 28899, 29146, 29393, 29640, 29887, 30134, 30381, 30628, 30875, 31122, 31369, 31616, 31863, 32110, 32357, 32604, 32851, 33098, 33345, 33592, 33839, 34086, 34333, 34580, 34827, 35074, 35321, 35568, 35815, 36062, 36309, 36556, 36803, 37050, 37297, 37544, 37791, 38038, 38285, 38532, 38779, 39026, 39273, 39520, 39767, 40014, 40261, 40508, 40755, 41002, 41249, 41496, 41743, 41990, 42237, 42484, 42731, 42978, 43225, 43472, 43719, 43966, 44213, 44460, 44707, 44954, 45201, 45448, 45695, 45942, 46189, 46436, 46683, 46930, 47177, 47424, 47671, 47918, 48165, 48412, 48659, 48906, 49153, 49400, 49647, 49894, 50141, 50388, 50635, 50882, 51129, 51376, 51623, 51870, 52117, 52364, 52611, 52858, 53105, 53352, 53599, 53846, 54093, 54340, 54587, 54834, 55081, 55328, 55575, 55822, 56069, 56316, 56563, 56810, 57057, 57304, 57551, 57798, 58045, 58292, 58539, 58786, 59033, 59280, 59527, 59774, 60021, 60268, 60515, 60762, 61009, 61256, 61503, 61750, 61997, 62244, 62491, 62738, 62985, 
0, 248, 496, 744, 992, 1240, 1488, 1736, 1984, 2232, 2480, 2728, 2976, 3224, 3472, 3720, 3968, 4216, 4464, 4712, 4960, 5208, 5456, 5704, 5952, 6200, 6448, 6696, 6944, 7192, 7440, 7688, 7936, 8184, 8432, 8680, 8928, 9176, 9424, 9672, 9920, 10168, 10416, 10664, 10912, 11160, 11408, 11656, 11904, 12152, 12400, 12648, 12896, 13144, 13392, 13640, 13888, 14136, 14384, 14632, 14880, 15128, 15376, 15624, 15872, 16120, 16368, 16616, 16864, 17112, 17360, 17608, 17856, 18104, 18352, 18600, 18848, 19096, 19344, 19592, 19840, 20088, 20336, 20584, 20832, 21080, 21328, 21576, 21824, 22072, 22320, 22568, 22816, 23064, 23312, 23560, 23808, 24056, 24304, 24552, 24800, 25048, 25296, 25544, 25792, 26040, 26288, 26536, 26784, 27032, 27280, 27528, 27776, 28024, 28272, 28520, 28768, 29016, 29264, 29512, 29760, 30008, 30256, 30504, 30752, 31000, 31248, 31496, 31744, 31992, 32240, 32488, 32736, 32984, 33232, 33480, 33728, 33976, 34224, 34472, 34720, 34968, 35216, 35464, 35712, 35960, 36208, 36456, 36704, 36952, 37200, 37448, 37696, 37944, 38192, 38440, 38688, 38936, 39184, 39432, 39680, 39928, 40176, 40424, 40672, 40920, 41168, 41416, 41664, 41912, 42160, 42408, 42656, 42904, 43152, 43400, 43648, 43896, 44144, 44392, 44640, 44888, 45136, 45384, 45632, 45880, 46128, 46376, 46624, 46872, 47120, 47368, 47616, 47864, 48112, 48360, 48608, 48856, 49104, 49352, 49600, 49848, 50096, 50344, 50592, 50840, 51088, 51336, 51584, 51832, 52080, 52328, 52576, 52824, 53072, 53320, 53568, 53816, 54064, 54312, 54560, 54808, 55056, 55304, 55552, 55800, 56048, 56296, 56544, 56792, 57040, 57288, 57536, 57784, 58032, 58280, 58528, 58776, 59024, 59272, 59520, 59768, 60016, 60264, 60512, 60760, 61008, 61256, 61504, 61752, 62000, 62248, 62496, 62744, 62992, 63240, 
0, 249, 498, 747, 996, 1245, 1494, 1743, 1992, 2241, 2490, 2739, 2988, 3237, 3486, 3735, 3984, 4233, 4482, 4731, 4980, 5229, 5478, 5727, 5976, 6225, 6474, 6723, 6972, 7221, 7470, 7719, 7968, 8217, 8466, 8715, 8964, 9213, 9462, 9711, 9960, 10209, 10458, 10707, 10956, 11205, 11454, 11703, 11952, 12201, 12450, 12699, 12948, 13197, 13446, 13695, 13944, 14193, 14442, 14691, 14940, 15189, 15438, 15687, 15936, 16185, 16434, 16683, 16932, 17181, 17430, 17679, 17928, 18177, 18426, 18675, 18924, 19173, 19422, 19671, 19920, 20169, 20418, 20667, 20916, 21165, 21414, 21663, 21912, 22161, 22410, 22659, 22908, 23157, 23406, 23655, 23904, 24153, 24402, 24651, 24900, 25149, 25398, 25647, 25896, 26145, 26394, 26643, 26892, 27141, 27390, 27639, 27888, 28137, 28386, 28635, 28884, 29133, 29382, 29631, 29880, 30129, 30378, 30627, 30876, 31125, 31374, 31623, 31872, 32121, 32370, 32619, 32868, 33117, 33366, 33615, 33864, 34113, 34362, 34611, 34860, 35109, 35358, 35607, 35856, 36105, 36354, 36603, 36852, 37101, 37350, 37599, 37848, 38097, 38346, 38595, 38844, 39093, 39342, 39591, 39840, 40089, 40338, 40587, 40836, 41085, 41334, 41583, 41832, 42081, 42330, 42579, 42828, 43077, 43326, 43575, 43824, 44073, 44322, 44571, 44820, 45069, 45318, 45567, 45816, 46065, 46314, 46563, 46812, 47061, 47310, 47559, 47808, 48057, 48306, 48555, 48804, 49053, 49302, 49551, 49800, 50049, 50298, 50547, 50796, 51045, 51294, 51543, 51792, 52041, 52290, 52539, 52788, 53037, 53286, 53535, 53784, 54033, 54282, 54531, 54780, 55029, 55278, 55527, 55776, 56025, 56274, 56523, 56772, 57021, 57270, 57519, 57768, 58017, 58266, 58515, 58764, 59013, 59262, 59511, 59760, 60009, 60258, 60507, 60756, 61005, 61254, 61503, 61752, 62001, 62250, 62499, 62748, 62997, 63246, 63495, 
0, 250, 500, 750, 1000, 1250, 1500, 1750, 2000, 2250, 2500, 2750, 3000, 3250, 3500, 3750, 4000, 4250, 4500, 4750, 5000, 5250, 5500, 5750, 6000, 6250, 6500, 6750, 7000, 7250, 7500, 7750, 8000, 8250, 8500, 8750, 9000, 9250, 9500, 9750, 10000, 10250, 10500, 10750, 11000, 11250, 11500, 11750, 12000, 12250, 12500, 12750, 13000, 13250, 13500, 13750, 14000, 14250, 14500, 14750, 15000, 15250, 15500, 15750, 16000, 16250, 16500, 16750, 17000, 17250, 17500, 17750, 18000, 18250, 18500, 18750, 19000, 19250, 19500, 19750, 20000, 20250, 20500, 20750, 21000, 21250, 21500, 21750, 22000, 22250, 22500, 22750, 23000, 23250, 23500, 23750, 24000, 24250, 24500, 24750, 25000, 25250, 25500, 25750, 26000, 26250, 26500, 26750, 27000, 27250, 27500, 27750, 28000, 28250, 28500, 28750, 29000, 29250, 29500, 29750, 30000, 30250, 30500, 30750, 31000, 31250, 31500, 31750, 32000, 32250, 32500, 32750, 33000, 33250, 33500, 33750, 34000, 34250, 34500, 34750, 35000, 35250, 35500, 35750, 36000, 36250, 36500, 36750, 37000, 37250, 37500, 37750, 38000, 38250, 38500, 38750, 39000, 39250, 39500, 39750, 40000, 40250, 40500, 40750, 41000, 41250, 41500, 41750, 42000, 42250, 42500, 42750, 43000, 43250, 43500, 43750, 44000, 44250, 44500, 44750, 45000, 45250, 45500, 45750, 46000, 46250, 46500, 46750, 47000, 47250, 47500, 47750, 48000, 48250, 48500, 48750, 49000, 49250, 49500, 49750, 50000, 50250, 50500, 50750, 51000, 51250, 51500, 51750, 52000, 52250, 52500, 52750, 53000, 53250, 53500, 53750, 54000, 54250, 54500, 54750, 55000, 55250, 55500, 55750, 56000, 56250, 56500, 56750, 57000, 57250, 57500, 57750, 58000, 58250, 58500, 58750, 59000, 59250, 59500, 59750, 60000, 60250, 60500, 60750, 61000, 61250, 61500, 61750, 62000, 62250, 62500, 62750, 63000, 63250, 63500, 63750, 
0, 251, 502, 753, 1004, 1255, 1506, 1757, 2008, 2259, 2510, 2761, 3012, 3263, 3514, 3765, 4016, 4267, 4518, 4769, 5020, 5271, 5522, 5773, 6024, 6275, 6526, 6777, 7028, 7279, 7530, 7781, 8032, 8283, 8534, 8785, 9036, 9287, 9538, 9789, 10040, 10291, 10542, 10793, 11044, 11295, 11546, 11797, 12048, 12299, 12550, 12801, 13052, 13303, 13554, 13805, 14056, 14307, 14558, 14809, 15060, 15311, 15562, 15813, 16064, 16315, 16566, 16817, 17068, 17319, 17570, 17821, 18072, 18323, 18574, 18825, 19076, 19327, 19578, 19829, 20080, 20331, 20582, 20833, 21084, 21335, 21586, 21837, 22088, 22339, 22590, 22841, 23092, 23343, 23594, 23845, 24096, 24347, 24598, 24849, 25100, 25351, 25602, 25853, 26104, 26355, 26606, 26857, 27108, 27359, 27610, 27861, 28112, 28363, 28614, 28865, 29116, 29367, 29618, 29869, 30120, 30371, 30622, 30873, 31124, 31375, 31626, 31877, 32128, 32379, 32630, 32881, 33132, 33383, 33634, 33885, 34136, 34387, 34638, 34889, 35140, 35391, 35642, 35893, 36144, 36395, 36646, 36897, 37148, 37399, 37650, 37901, 38152, 38403, 38654, 38905, 39156, 39407, 39658, 39909, 40160, 40411, 40662, 40913, 41164, 41415, 41666, 41917, 42168, 42419, 42670, 42921, 43172, 43423, 43674, 43925, 44176, 44427, 44678, 44929, 45180, 45431, 45682, 45933, 46184, 46435, 46686, 46937, 47188, 47439, 47690, 47941, 48192, 48443, 48694, 48945, 49196, 49447, 49698, 49949, 50200, 50451, 50702, 50953, 51204, 51455, 51706, 51957, 52208, 52459, 52710, 52961, 53212, 53463, 53714, 53965, 54216, 54467, 54718, 54969, 55220, 55471, 55722, 55973, 56224, 56475, 56726, 56977, 57228, 57479, 57730, 57981, 58232, 58483, 58734, 58985, 59236, 59487, 59738, 59989, 60240, 60491, 60742, 60993, 61244, 61495, 61746, 61997, 62248, 62499, 62750, 63001, 63252, 63503, 63754, 64005, 
0, 252, 504, 756, 1008, 1260, 1512, 1764, 2016, 2268, 2520, 2772, 3024, 3276, 3528, 3780, 4032, 4284, 4536, 4788, 5040, 5292, 5544, 5796, 6048, 6300, 6552, 6804, 7056, 7308, 7560, 7812, 8064, 8316, 8568, 8820, 9072, 9324, 9576, 9828, 10080, 10332, 10584, 10836, 11088, 11340, 11592, 11844, 12096, 12348, 12600, 12852, 13104, 13356, 13608, 13860, 14112, 14364, 14616, 14868, 15120, 15372, 15624, 15876, 16128, 16380, 16632, 16884, 17136, 17388, 17640, 17892, 18144, 18396, 18648, 18900, 19152, 19404, 19656, 19908, 20160, 20412, 20664, 20916, 21168, 21420, 21672, 21924, 22176, 22428, 22680, 22932, 23184, 23436, 23688, 23940, 24192, 24444, 24696, 24948, 25200, 25452, 25704, 25956, 26208, 26460, 26712, 26964, 27216, 27468, 27720, 27972, 28224, 28476, 28728, 28980, 29232, 29484, 29736, 29988, 30240, 30492, 30744, 30996, 31248, 31500, 31752, 32004, 32256, 32508, 32760, 33012, 33264, 33516, 33768, 34020, 34272, 34524, 34776, 35028, 35280, 35532, 35784, 36036, 36288, 36540, 36792, 37044, 37296, 37548, 37800, 38052, 38304, 38556, 38808, 39060, 39312, 39564, 39816, 40068, 40320, 40572, 40824, 41076, 41328, 41580, 41832, 42084, 42336, 42588, 42840, 43092, 43344, 43596, 43848, 44100, 44352, 44604, 44856, 45108, 45360, 45612, 45864, 46116, 46368, 46620, 46872, 47124, 47376, 47628, 47880, 48132, 48384, 48636, 48888, 49140, 49392, 49644, 49896, 50148, 50400, 50652, 50904, 51156, 51408, 51660, 51912, 52164, 52416, 52668, 52920, 53172, 53424, 53676, 53928, 54180, 54432, 54684, 54936, 55188, 55440, 55692, 55944, 56196, 56448, 56700, 56952, 57204, 57456, 57708, 57960, 58212, 58464, 58716, 58968, 59220, 59472, 59724, 59976, 60228, 60480, 60732, 60984, 61236, 61488, 61740, 61992, 62244, 62496, 62748, 63000, 63252, 63504, 63756, 64008, 64260, 
0, 253, 506, 759, 1012, 1265, 1518, 1771, 2024, 2277, 2530, 2783, 3036, 3289, 3542, 3795, 4048, 4301, 4554, 4807, 5060, 5313, 5566, 5819, 6072, 6325, 6578, 6831, 7084, 7337, 7590, 7843, 8096, 8349, 8602, 8855, 9108, 9361, 9614, 9867, 10120, 10373, 10626, 10879, 11132, 11385, 11638, 11891, 12144, 12397, 12650, 12903, 13156, 13409, 13662, 13915, 14168, 14421, 14674, 14927, 15180, 15433, 15686, 15939, 16192, 16445, 16698, 16951, 17204, 17457, 17710, 17963, 18216, 18469, 18722, 18975, 19228, 19481, 19734, 19987, 20240, 20493, 20746, 20999, 21252, 21505, 21758, 22011, 22264, 22517, 22770, 23023, 23276, 23529, 23782, 24035, 24288, 24541, 24794, 25047, 25300, 25553, 25806, 26059, 26312, 26565, 26818, 27071, 27324, 27577, 27830, 28083, 28336, 28589, 28842, 29095, 29348, 29601, 29854, 30107, 30360, 30613, 30866, 31119, 31372, 31625, 31878, 32131, 32384, 32637, 32890, 33143, 33396, 33649, 33902, 34155, 34408, 34661, 34914, 35167, 35420, 35673, 35926, 36179, 36432, 36685, 36938, 37191, 37444, 37697, 37950, 38203, 38456, 38709, 38962, 39215, 39468, 39721, 39974, 40227, 40480, 40733, 40986, 41239, 41492, 41745, 41998, 42251, 42504, 42757, 43010, 43263, 43516, 43769, 44022, 44275, 44528, 44781, 45034, 45287, 45540, 45793, 46046, 46299, 46552, 46805, 47058, 47311, 47564, 47817, 48070, 48323, 48576, 48829, 49082, 49335, 49588, 49841, 50094, 50347, 50600, 50853, 51106, 51359, 51612, 51865, 52118, 52371, 52624, 52877, 53130, 53383, 53636, 53889, 54142, 54395, 54648, 54901, 55154, 55407, 55660, 55913, 56166, 56419, 56672, 56925, 57178, 57431, 57684, 57937, 58190, 58443, 58696, 58949, 59202, 59455, 59708, 59961, 60214, 60467, 60720, 60973, 61226, 61479, 61732, 61985, 62238, 62491, 62744, 62997, 63250, 63503, 63756, 64009, 64262, 64515, 
0, 254, 508, 762, 1016, 1270, 1524, 1778, 2032, 2286, 2540, 2794, 3048, 3302, 3556, 3810, 4064, 4318, 4572, 4826, 5080, 5334, 5588, 5842, 6096, 6350, 6604, 6858, 7112, 7366, 7620, 7874, 8128, 8382, 8636, 8890, 9144, 9398, 9652, 9906, 10160, 10414, 10668, 10922, 11176, 11430, 11684, 11938, 12192, 12446, 12700, 12954, 13208, 13462, 13716, 13970, 14224, 14478, 14732, 14986, 15240, 15494, 15748, 16002, 16256, 16510, 16764, 17018, 17272, 17526, 17780, 18034, 18288, 18542, 18796, 19050, 19304, 19558, 19812, 20066, 20320, 20574, 20828, 21082, 21336, 21590, 21844, 22098, 22352, 22606, 22860, 23114, 23368, 23622, 23876, 24130, 24384, 24638, 24892, 25146, 25400, 25654, 25908, 26162, 26416, 26670, 26924, 27178, 27432, 27686, 27940, 28194, 28448, 28702, 28956, 29210, 29464, 29718, 29972, 30226, 30480, 30734, 30988, 31242, 31496, 31750, 32004, 32258, 32512, 32766, 33020, 33274, 33528, 33782, 34036, 34290, 34544, 34798, 35052, 35306, 35560, 35814, 36068, 36322, 36576, 36830, 37084, 37338, 37592, 37846, 38100, 38354, 38608, 38862, 39116, 39370, 39624, 39878, 40132, 40386, 40640, 40894, 41148, 41402, 41656, 41910, 42164, 42418, 42672, 42926, 43180, 43434, 43688, 43942, 44196, 44450, 44704, 44958, 45212, 45466, 45720, 45974, 46228, 46482, 46736, 46990, 47244, 47498, 47752, 48006, 48260, 48514, 48768, 49022, 49276, 49530, 49784, 50038, 50292, 50546, 50800, 51054, 51308, 51562, 51816, 52070, 52324, 52578, 52832, 53086, 53340, 53594, 53848, 54102, 54356, 54610, 54864, 55118, 55372, 55626, 55880, 56134, 56388, 56642, 56896, 57150, 57404, 57658, 57912, 58166, 58420, 58674, 58928, 59182, 59436, 59690, 59944, 60198, 60452, 60706, 60960, 61214, 61468, 61722, 61976, 62230, 62484, 62738, 62992, 63246, 63500, 63754, 64008, 64262, 64516, 64770, 
0, 255, 510, 765, 1020, 1275, 1530, 1785, 2040, 2295, 2550, 2805, 3060, 3315, 3570, 3825, 4080, 4335, 4590, 4845, 5100, 5355, 5610, 5865, 6120, 6375, 6630, 6885, 7140, 7395, 7650, 7905, 8160, 8415, 8670, 8925, 9180, 9435, 9690, 9945, 10200, 10455, 10710, 10965, 11220, 11475, 11730, 11985, 12240, 12495, 12750, 13005, 13260, 13515, 13770, 14025, 14280, 14535, 14790, 15045, 15300, 15555, 15810, 16065, 16320, 16575, 16830, 17085, 17340, 17595, 17850, 18105, 18360, 18615, 18870, 19125, 19380, 19635, 19890, 20145, 20400, 20655, 20910, 21165, 21420, 21675, 21930, 22185, 22440, 22695, 22950, 23205, 23460, 23715, 23970, 24225, 24480, 24735, 24990, 25245, 25500, 25755, 26010, 26265, 26520, 26775, 27030, 27285, 27540, 27795, 28050, 28305, 28560, 28815, 29070, 29325, 29580, 29835, 30090, 30345, 30600, 30855, 31110, 31365, 31620, 31875, 32130, 32385, 32640, 32895, 33150, 33405, 33660, 33915, 34170, 34425, 34680, 34935, 35190, 35445, 35700, 35955, 36210, 36465, 36720, 36975, 37230, 37485, 37740, 37995, 38250, 38505, 38760, 39015, 39270, 39525, 39780, 40035, 40290, 40545, 40800, 41055, 41310, 41565, 41820, 42075, 42330, 42585, 42840, 43095, 43350, 43605, 43860, 44115, 44370, 44625, 44880, 45135, 45390, 45645, 45900, 46155, 46410, 46665, 46920, 47175, 47430, 47685, 47940, 48195, 48450, 48705, 48960, 49215, 49470, 49725, 49980, 50235, 50490, 50745, 51000, 51255, 51510, 51765, 52020, 52275, 52530, 52785, 53040, 53295, 53550, 53805, 54060, 54315, 54570, 54825, 55080, 55335, 55590, 55845, 56100, 56355, 56610, 56865, 57120, 57375, 57630, 57885, 58140, 58395, 58650, 58905, 59160, 59415, 59670, 59925, 60180, 60435, 60690, 60945, 61200, 61455, 61710, 61965, 62220, 62475, 62730, 62985, 63240, 63495, 63750, 64005, 64260, 64515, 64770, 65025 );
 
BEGIN
 
	-- Instantiate the Unit Under Test (UUT)
   uut: entity work.hw_mul_pipelined 
   GENERIC MAP(
		  N => 8,
		  M => 8 )
   PORT MAP (
          rst => reset,
          clk => clk,
          validin => valid_in,
          a => a,
          b => b,
          validout => valid_out,
          q => q
        );

	stim_process: process
	begin
		reset <= '1';
		
		wait for 100 ns;
		
		reset <= '0';
   
		for I in 0 to 255 loop
			for J in 0 to 255 loop
				clk <= '0';
				valid_in <= '1';
				a <= to_unsigned(I, 8);
				b <= to_unsigned(J, 8);
				wait for clk_period/2;
				clk <= '1';
				wait for clk_period/2;
			end loop;
		end loop;
		
		valid_in <= '0';
		
		for J in 0 to 15 loop
			clk <= '0';
			wait for clk_period/2;
			clk <= '1';
			wait for clk_period/2;
		end loop;

		wait;
		
	end process stim_process;
   
	process(clk)
	begin
		if( falling_edge( clk ) ) then
			if( valid_out = '1' ) then
			
				assert q = to_unsigned(results(counter), 16)
					report "Wrong value. Expecting " & 
						integer'image(results(counter)) & 
						" is " & 
						integer'image(to_integer(q))
					severity warning;
					
				counter <= counter + 1;
			end if;
		end if;
	end process;

END;
