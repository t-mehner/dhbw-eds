----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 		Torben Mehner
-- 
-- Create Date:		07:40:50 10/02/2019 
-- Design Name:
-- Module Name:		led_out - Behavioral 
-- Project Name: 	01_led_out
-- Target Devices: 
-- Tool versions: 
-- Description: 
--
-- Dependencies: 
--
-- Revision: 
-- Revision 0.01 - File Created
-- Additional Comments: 
--
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx primitives in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity led_out is
    Port ( SW  : in  STD_LOGIC_VECTOR (7 downto 0);
           LED : out  STD_LOGIC_VECTOR (7 downto 0));
end led_out;

architecture Behavioral of led_out is

begin

	-- add logic statements here

end Behavioral;

